// Verilog
// c2670
// N in 233
// N out 140
// NtotalGates 1269

module c2670 (clk, en, N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, N37, N40, N43, N44,
			  N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76, N77, N78, N79, N80, 
			  N81, N82, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N111, N112, N113, N114,
			  N115, N116, N117, N118, N119, N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N138, N139, N140, N141, N142, N219, 
			  N224, N227, N230, N231, N234, N237, N241, N246, N253, N256, N259, N262, N263, N266, N269, N272, N275, N278, N281, N284, N287, N290, N294, N297, N301, 
			  N305, N309, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N143_I, N144_I, N145_I, N146_I, N147_I, N148_I, 
			  N149_I, N150_I, N151_I, N152_I, N153_I, N154_I, N155_I, N156_I, N157_I, N158_I, N159_I, N160_I, N161_I, N162_I, N163_I, N164_I, N165_I, N166_I, N167_I,
			  N168_I, N169_I, N170_I, N171_I, N172_I, N173_I, N174_I, N175_I, N176_I, N177_I, N178_I, N179_I, N180_I, N181_I, N182_I, N183_I, N184_I, N185_I, N186_I, N187_I, N188_I, N189_I, N190_I, N191_I, N192_I, N193_I, N194_I, N195_I, N196_I, N197_I, N198_I, N199_I, N200_I, N201_I, N202_I, N203_I, N204_I, N205_I, N206_I, N207_I, N208_I, N209_I, N210_I, N211_I, N212_I, N213_I, N214_I, N215_I, N216_I, N217_I, N218_I, N398, N400, N401, N419, N420, N456, N457, 
			  N458, N487, N488, N489, N490, N491, N492, N493, N494, N792, N799, N805, N1026, N1028, N1029, N1269, N1277, N1448, N1726, N1816, N1817, N1818, N1819, 
			  N1820, N1821, N1969, N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022, N2387, N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925, 
			  N2970, N2971, N3038, N3079, N3546, N3671, N3803, N3804, N3809, N3851, N3875, N3881, N3882, N143_O, N144_O, N145_O, N146_O, N147_O, N148_O, N149_O, 
			  N150_O, N151_O, N152_O, N153_O, N154_O, N155_O, N156_O, N157_O, N158_O, N159_O, N160_O, N161_O, N162_O, N163_O, N164_O, N165_O, N166_O, N167_O, N168_O,
			  N169_O, N170_O, N171_O, N172_O, N173_O, N174_O, N175_O, N176_O, N177_O, N178_O, N179_O, N180_O, N181_O, N182_O, N183_O, N184_O, N185_O, N186_O, N187_O,
			  N188_O, N189_O, N190_O, N191_O, N192_O, N193_O, N194_O, N195_O, N196_O, N197_O, N198_O, N199_O, N200_O, N201_O, N202_O, N203_O, N204_O, N205_O, N206_O,
			  N207_O, N208_O, N209_O, N210_O, N211_O, N212_O, N213_O, N214_O, N215_O, N216_O, N217_O, N218_O);

input clk, en, N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22, N23, N24, N25, N26,  N27, N28, N29, N32, N33, N34, N35, N36, N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54,  N55, N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76, N77, N78,  N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N99, N100, N101, N102,  N103, N104, N105, N106, N107, N108, N111, N112, N113, N114,  N115, N116, N117, N118, N119, N120, N123, N124, N125, N126,  N127, N128, N129, N130, N131, N132, N135, N136, N137, N138,  N139, N140, N141, N142, N219, N224, N227, N230, N231, N234,  N237, N241, N246, N253, N256, N259, N262, N263, N266, N269,  N272, N275, N278, N281, N284, N287, N290, N294, N297, N301,  N305, N309, N313, N316, N319, N322, N325, N328, N331, N334,  N337, N340, N343, N346, N349, N352, N355, N143_I, N144_I, N145_I,  N146_I, N147_I, N148_I, N149_I, N150_I, N151_I, N152_I, N153_I, N154_I, N155_I,  N156_I, N157_I, N158_I, N159_I, N160_I, N161_I, N162_I, N163_I, N164_I, N165_I,  N166_I, N167_I, N168_I, N169_I, N170_I, N171_I, N172_I, N173_I, N174_I, N175_I,  N176_I, N177_I, N178_I, N179_I, N180_I, N181_I, N182_I, N183_I, N184_I, N185_I,  N186_I, N187_I, N188_I, N189_I, N190_I, N191_I, N192_I, N193_I, N194_I, N195_I,  N196_I, N197_I, N198_I, N199_I, N200_I, N201_I, N202_I, N203_I, N204_I, N205_I,  N206_I, N207_I, N208_I, N209_I, N210_I, N211_I, N212_I, N213_I, N214_I, N215_I,  N216_I, N217_I, N218_I; 

output N398, N400, N401, N419, N420, N456, N457, N458, N487, N488, N489, N490, N491, N492, N493, N494, N792, N799, N805, N1026, N1028, N1029, N1269, N1277, N1448, N1726, N1816, N1817, N1818, N1819, N1820, N1821, N1969, N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022, N2387, N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925, N2970, N2971, N3038, N3079, N3546, N3671, N3803, N3804, N3809, N3851, N3875, N3881, N3882, N143_O, N144_O, N145_O, N146_O, N147_O, N148_O, N149_O, N150_O, N151_O, N152_O, N153_O, N154_O, N155_O, N156_O, N157_O, N158_O, N159_O, N160_O, N161_O, N162_O, N163_O, N164_O, N165_O, N166_O, N167_O, N168_O, N169_O, N170_O, N171_O, N172_O, N173_O, N174_O, N175_O, N176_O, N177_O, N178_O, N179_O, N180_O, N181_O, N182_O, N183_O, N184_O, N185_O, N186_O, N187_O, N188_O, N189_O, N190_O, N191_O, N192_O, N193_O, N194_O, N195_O, N196_O, N197_O, N198_O, N199_O, N200_O, N201_O, N202_O, N203_O, N204_O, N205_O, N206_O, N207_O, N208_O, N209_O, N210_O, N211_O, N212_O, N213_O, N214_O, N215_O, N216_O, N217_O, N218_O;

wire N1880, N2880, error, dN1, dN2, dN3, dN4, dN5, dN6, dN7, dN8, dN11, dN14, dN15, dN16, dN19, dN20, dN21, dN22, dN23, dN24, dN25, dN26,  dN27, dN28, dN29, dN32, dN33, dN34, dN35, dN36, dN37, dN40, dN43, dN44, dN47, dN48, dN49, dN50, dN51, dN52, dN53, dN54,  dN55, dN56, dN57, dN60, dN61, dN62, dN63, dN64, dN65, dN66, dN67, dN68, dN69, dN72, dN73, dN74, dN75, dN76, dN77, dN78,  dN79, dN80, dN81, dN82, dN85, dN86, dN87, dN88, dN89, dN90, dN91, dN92, dN93, dN94, dN95, dN96, dN99, dN100, dN101, dN102,  dN103, dN104, dN105, dN106, dN107, dN108, dN111, dN112, dN113, dN114,  dN115, dN116, dN117, dN118, dN119, dN120, dN123, dN124, dN125, dN126,  dN127, dN128, dN129, dN130, dN131, dN132, dN135, dN136, dN137, dN138,  dN139, dN140, dN141, dN142, dN219, dN224, dN227, dN230, dN231, dN234,  dN237, dN241, dN246, dN253, dN256, dN259, dN262, dN263, dN266, dN269,  dN272, dN275, dN278, dN281, dN284, dN287, dN290, dN294, dN297, dN301,  dN305, dN309, dN313, dN316, dN319, dN322, dN325, dN328, dN331, dN334,  dN337, dN340, dN343, dN346, dN349, dN352, dN355, dN143_I, dN144_I, dN145_I,  dN146_I, dN147_I, dN148_I, dN149_I, dN150_I, dN151_I, dN152_I, dN153_I, dN154_I, dN155_I,  dN156_I, dN157_I, dN158_I, dN159_I, dN160_I, dN161_I, dN162_I, dN163_I, dN164_I, dN165_I,  dN166_I, dN167_I, dN168_I, dN169_I, dN170_I, dN171_I, dN172_I, dN173_I, dN174_I, dN175_I,  dN176_I, dN177_I, dN178_I, dN179_I, dN180_I, dN181_I, dN182_I, dN183_I, dN184_I, dN185_I,  dN186_I, dN187_I, dN188_I, dN189_I, dN190_I, dN191_I, dN192_I, dN193_I, dN194_I, dN195_I,  dN196_I, dN197_I, dN198_I, dN199_I, dN200_I, dN201_I, dN202_I, dN203_I, dN204_I, dN205_I,  dN206_I, dN207_I, dN208_I, dN209_I, dN210_I, dN211_I, dN212_I, dN213_I, dN214_I, dN215_I,  dN216_I, dN217_I, dN218_I, dN398, dN400, dN401, dN419, dN420, dN456, dN457, dN458, dN487, dN488, dN489, dN490, dN491, dN492, dN493, dN494, dN792, dN799, dN805, dN1026, dN1028, dN1029, dN1269, dN1277, dN1448, dN1726, dN1816, dN1817, dN1818, dN1819, dN1820, dN1821, dN1969, dN1970, dN1971, dN2010, dN2012, dN2014, dN2016, dN2018, dN2020, dN2022, dN2387, dN2388, dN2389, dN2390, dN2496, dN2643, dN2644, dN2891, dN2925, dN2970, dN2971, dN3038, dN3079, dN3546, dN3671, dN3803, dN3804, dN3809, dN3851, dN3875, dN3881, dN3882, dN143_O, dN144_O, dN145_O, dN146_O, dN147_O, dN148_O, dN149_O, dN150_O, dN151_O, dN152_O, dN153_O, dN154_O, dN155_O, dN156_O, dN157_O, dN158_O, dN159_O, dN160_O, dN161_O, dN162_O, dN163_O, dN164_O, dN165_O, dN166_O, dN167_O, dN168_O, dN169_O, dN170_O, dN171_O, dN172_O, dN173_O, dN174_O, dN175_O, dN176_O, dN177_O, dN178_O, dN179_O, dN180_O, dN181_O, dN182_O, dN183_O, dN184_O, dN185_O, dN186_O, dN187_O, dN188_O, dN189_O, dN190_O, dN191_O, dN192_O, dN193_O, dN194_O, dN195_O, dN196_O, dN197_O, dN198_O, dN199_O, dN200_O, dN201_O, dN202_O, dN203_O, dN204_O, dN205_O, dN206_O, dN207_O, dN208_O, dN209_O, dN210_O, dN211_O, dN212_O, dN213_O, dN214_O, dN215_O, dN216_O, dN217_O, dN218_O, N405, N408, N425, N485, N486, N495, N496, N499, N500, N503, N506, N509, N521, N533, N537, N543, N544, N547, N550, N562, N574, N578, N582, N594, N606, N607, N608, N609, N610, N611, N612, N613, N625, N637, N643, N650, N651, N655, N659, N663, N667, N671, N675, N679, N683, N687, N693, N699, N705, N711, N715, N719, N723, N727, N730, N733, N734, N735, N738, N741, N744, N747, N750, N753, N756, N759, N762, N765, N768, N771, N774, N777, N780, N783, N786, N800, N900, N901, N902, N903, N904, N905, N998, N999, N1027, N1032, N1033, N1034, N1037, N1042, N1053, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1075, N1086, N1097, N1098, N1099, N1100, N1101, N1102, N1113, N1124, N1125, N1126, N1127, N1128, N1129, N1133, N1137, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1157, N1168, N1169, N1170, N1171, N1172, N1173, N1178, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1195, N1200, N1205, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1219, N1222, N1225, N1228, N1231, N1234, N1237, N1240, N1243, N1246, N1249, N1250, N1251, N1254, N1257, N1260, N1263, N1266, N1275, N1276, N1302, N1351, N1352, N1353, N1354, N1355, N1395, N1396, N1397, N1398, N1399, N1422, N1423, N1424, N1425, N1426, N1427, N1440, N1441, N1449, N1450, N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462, N1463, N1464, N1465, N1466, N1467, N1468, N1469, N1470, N1471, N1472, N1473, N1474, N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483, N1484, N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493, N1494, N1495, N1496, N1499, N1502, N1506, N1510, N1513, N1516, N1519, N1520, N1521, N1522, N1523, N1524, N1525, N1526, N1527, N1528, N1529, N1530, N1531, N1532, N1533, N1534, N1535, N1536, N1537, N1538, N1539, N1540, N1541, N1542, N1543, N1544, N1545, N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1553, N1557, N1561, N1564, N1565, N1566, N1567, N1568, N1569, N1570, N1571, N1572, N1573, N1574, N1575, N1576, N1577, N1578, N1581, N1582, N1585, N1588, N1591, N1596, N1600, N1606, N1612, N1615, N1619, N1624, N1628, N1631, N1634, N1637, N1642, N1647, N1651, N1656, N1676, N1681, N1686, N1690, N1708, N1770, N1773, N1776, N1777, N1778, N1781, N1784, N1785, N1795, N1798, N1801, N1804, N1807, N1808, N1809, N1810, N1811, N1813, N1814, N1815, N1822, N1823, N1824, N1827, N1830, N1831, N1832, N1833, N1836, N1841, N1848, N1852, N1856, N1863, N1870, N1875, N12670, N1885, N1888, N1891, N1894, N1897, N1908, N1909, N1910, N1911, N1912, N1913, N1914, N1915, N1916, N1917, N1918, N1919, N1928, N1929, N1930, N1931, N1932, N1933, N1934, N1935, N1936, N1939, N1940, N1941, N1942, N1945, N1948, N1951, N1954, N1957, N1960, N1963, N1966, N2028, N2029, N2030, N2031, N2032, N2033, N2034, N2040, N2041, N2042, N2043, N2046, N2049, N2052, N2055, N2058, N2061, N2064, N2067, N2070, N2073, N2076, N2079, N2095, N2098, N2101, N2104, N2107, N2110, N2113, N2119, N2120, N2125, N2126, N2127, N2128, N2135, N2141, N2144, N2147, N2150, N2153, N2154, N2155, N2156, N2157, N2158, N2171, N2172, N2173, N2174, N2175, N2176, N2177, N2178, N2185, N2188, N2191, N2194, N2197, N2200, N2201, N2204, N2207, N2210, N2213, N2216, N2219, N2234, N2235, N2236, N2237, N2250, N2266, N2269, N2291, N2294, N2297, N2298, N2300, N2301, N2302, N2303, N2304, N2305, N2306, N2307, N2308, N2309, N2310, N2311, N2312, N2313, N2314, N2315, N2316, N2317, N2318, N2319, N2320, N2321, N2322, N2323, N2324, N2325, N2326, N2327, N2328, N2329, N2330, N2331, N2332, N2333, N2334, N2335, N2336, N2337, N2338, N2339, N2340, N2354, N2355, N2356, N2357, N2358, N2359, N2364, N2365, N2366, N2367, N2368, N2372, N2373, N2374, N2375, N2376, N2377, N2382, N2386, N2391, N2395, N2400, N2403, N2406, N2407, N2408, N2409, N2410, N2411, N2412, N2413, N2414, N2415, N2416, N2417, N2421, N2425, N2428, N2429, N2430, N2431, N2432, N2433, N2434, N2437, N2440, N2443, N2446, N2449, N2452, N2453, N2454, N2457, N2460, N2463, N2466, N2469, N2472, N2475, N2478, N2481, N2484, N2487, N2490, N2493, N2503, N2504, N2510, N2511, N2521, N2528, N2531, N2534, N2537, N2540, N2544, N2545, N2546, N2547, N2548, N2549, N2550, N2551, N2552, N2553, N2563, N2564, N2565, N2566, N2567, N2568, N2579, N2603, N2607, N2608, N2609, N2610, N2611, N2612, N2613, N2617, N2618, N2619, N2620, N2621, N2624, N2628, N2629, N2630, N2631, N2632, N2633, N2634, N2635, N2636, N2638, N2645, N2646, N2652, N2655, N2656, N2659, N2663, N2664, N2665, N2666, N2667, N2668, N2669, N2670, N2671, N2672, N2673, N2674, N2675, N2676, N2677, N2678, N2679, N2680, N2681, N2684, N2687, N2690, N2693, N2694, N2695, N2696, N2697, N2698, N2699, N2700, N2701, N2702, N2703, N2706, N2707, N2708, N2709, N2710, N2719, N2720, N2726, N2729, N2738, N2743, N2747, N2748, N2749, N2750, N2751, N2760, N2761, N2766, N2771, N2772, N2773, N2774, N2775, N2776, N2777, N2778, N2781, N2782, N2783, N2784, N2789, N2790, N2791, N2792, N2793, N2796, N2800, N2803, N2806, N2809, N2810, N2811, N2812, N2817, N2820, N2826, N2829, N2830, N2831, N2837, N2838, N2839, N2840, N2841, N2844, N2854, N2859, N2869, N2874, N2877, N22670, N2881, N2882, N2885, N2888, N2894, N2895, N2896, N2897, N2898, N2899, N2900, N2901, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2931, N2938, N2939, N2963, N2972, N2975, N2978, N2981, N2984, N2985, N2986, N2989, N2992, N2995, N2998, N3001, N3004, N3007, N3008, N3009, N3010, N3013, N3016, N3019, N3022, N3025, N3028, N3029, N3030, N3035, N3036, N3037, N3039, N3044, N3045, N3046, N3047, N3048, N3049, N3050, N3053, N3054, N3055, N3056, N3057, N3058, N3059, N3060, N3061, N3064, N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, N3075, N3076, N3088, N3091, N3110, N3113, N3137, N3140, N3143, N3146, N3149, N3152, N3157, N3160, N3163, N3166, N3169, N3172, N3175, N3176, N3177, N3178, N3180, N3187, N3188, N3189, N3190, N3191, N3192, N3193, N3194, N3195, N3196, N3197, N3208, N3215, N3216, N3217, N3218, N3219, N3220, N3222, N3223, N3230, N3231, N3238, N3241, N3244, N3247, N3250, N3253, N3256, N3259, N3262, N3265, N3268, N3271, N3274, N3277, N3281, N3282, N3283, N3284, N3286, N3288, N3289, N3291, N3293, N3295, N3296, N3299, N3301, N3302, N3304, N3306, N3308, N3309, N3312, N3314, N3315, N3318, N3321, N3324, N3327, N3330, N3333, N3334, N3335, N3336, N3337, N3340, N3344, N3348, N3352, N3356, N3360, N3364, N3367, N3370, N3374, N3378, N3382, N3386, N3390, N3394, N3397, N3400, N3401, N3402, N3403, N3404, N3405, N3406, N3409, N3410, N3412, N3414, N3416, N3418, N3420, N3422, N3428, N3430, N3432, N3434, N3436, N3438, N3440, N3450, N3453, N3456, N3459, N3478, N3479, N3480, N3481, N3482, N3483, N3484, N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, N3493, N3494, N3496, N3498, N3499, N3500, N3501, N3502, N3503, N3504, N3505, N3506, N3507, N3508, N3509, N3510, N3511, N3512, N3513, N3515, N3517, N3522, N3525, N3528, N3531, N3534, N3537, N3540, N3543, N3551, N3552, N3553, N3554, N3555, N3556, N3557, N3558, N3559, N3563, N3564, N3565, N3566, N3567, N3568, N3569, N3570, N3576, N3579, N3585, N3588, N3592, N3593, N3594, N3595, N3596, N3597, N3598, N3599, N3600, N3603, N3608, N3612, N3615, N3616, N3622, N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3640, N3644, N3647, N3648, N3654, N3661, N3662, N3667, N3668, N3669, N3670, N3691, N3692, N3693, N3694, N3695, N3696, N3697, N3716, N3717, N3718, N3719, N3720, N3721, N3722, N3723, N3726, N3727, N3728, N3729, N3730, N3731, N3732, N3733, N3734, N3735, N3736, N3737, N3740, N3741, N3742, N3743, N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3753, N3754, N3758, N3761, N3762, N3767, N3771, N3774, N3775, N3778, N3779, N3780, N3790, N3793, N3794, N3802, N3805, N3806, N3807, N3808, N3811, N3812, N3813, N3814, N3815, N3816, N3817, N3818, N3819, N3820, N3821, N3822, N3823, N3826, N3827, N3834, N3835, N3836, N3837, N3838, N3839, N3840, N3843, N3852, N3857, N3858, N3859, N3864, N3869, N3870, N3876, N3877;

buf BUFF1_1 (dN398, dN219);
buf BUFF1_2 (dN400, dN219);
buf BUFF1_3 (dN401, dN219);
and AND2_4 (N405, dN1, dN3);
not NOT1_5 (N408, dN230);
buf BUFF1_6 (dN419, dN253);
buf BUFF1_7 (dN420, dN253);
not NOT1_8 (N425, dN262);
buf BUFF1_9 (dN456, dN290);
buf BUFF1_10 (dN457, dN290);
buf BUFF1_11 (dN458, dN290);
and AND4_12 (N485, dN309, dN305, dN301, dN297);
not NOT1_13 (N486, N405);
not NOT1_14 (dN487, dN44);
not NOT1_15 (dN488, dN132);
not NOT1_16 (dN489, dN82);
not NOT1_17 (dN490, dN96);
not NOT1_18 (dN491, dN69);
not NOT1_19 (dN492, dN120);
not NOT1_20 (dN493, dN57);
not NOT1_21 (dN494, dN108);
and AND3_22 (N495, dN2, dN15, dN237);
buf BUFF1_23 (N496, dN237);
and AND2_24 (N499, dN37, dN37);
buf BUFF1_25 (N500, dN219);
buf BUFF1_26 (N503, dN8);
buf BUFF1_27 (N506, dN8);
buf BUFF1_28 (N509, dN227);
buf BUFF1_29 (N521, dN234);
not NOT1_30 (N533, dN241);
not NOT1_31 (N537, dN246);
and AND2_32 (N543, dN11, dN246);
and AND4_33 (N544, dN132, dN82, dN96, dN44);
and AND4_34 (N547, dN120, dN57, dN108, dN69);
buf BUFF1_35 (N550, dN227);
buf BUFF1_36 (N562, dN234);
not NOT1_37 (N574, dN256);
not NOT1_38 (N578, dN259);
buf BUFF1_39 (N582, dN319);
buf BUFF1_40 (N594, dN322);
not NOT1_41 (N606, dN328);
not NOT1_42 (N607, dN331);
not NOT1_43 (N608, dN334);
not NOT1_44 (N609, dN337);
not NOT1_45 (N610, dN340);
not NOT1_46 (N611, dN343);
not NOT1_47 (N612, dN352);
buf BUFF1_48 (N613, dN319);
buf BUFF1_49 (N625, dN322);
buf BUFF1_50 (N637, dN16);
buf BUFF1_51 (N643, dN16);
not NOT1_52 (N650, dN355);
and AND2_53 (N651, dN7, dN237);
not NOT1_54 (N655, dN263);
not NOT1_55 (N659, dN266);
not NOT1_56 (N663, dN269);
not NOT1_57 (N667, dN272);
not NOT1_58 (N671, dN275);
not NOT1_59 (N675, dN278);
not NOT1_60 (N679, dN281);
not NOT1_61 (N683, dN284);
not NOT1_62 (N687, dN287);
buf BUFF1_63 (N693, dN29);
buf BUFF1_64 (N699, dN29);
not NOT1_65 (N705, dN294);
not NOT1_66 (N711, dN297);
not NOT1_67 (N715, dN301);
not NOT1_68 (N719, dN305);
not NOT1_69 (N723, dN309);
not NOT1_70 (N727, dN313);
not NOT1_71 (N730, dN316);
not NOT1_72 (N733, dN346);
not NOT1_73 (N734, dN349);
buf BUFF1_74 (N735, dN259);
buf BUFF1_75 (N738, dN256);
buf BUFF1_76 (N741, dN263);
buf BUFF1_77 (N744, dN269);
buf BUFF1_78 (N747, dN266);
buf BUFF1_79 (N750, dN275);
buf BUFF1_80 (N753, dN272);
buf BUFF1_81 (N756, dN281);
buf BUFF1_82 (N759, dN278);
buf BUFF1_83 (N762, dN287);
buf BUFF1_84 (N765, dN284);
buf BUFF1_85 (N768, dN294);
buf BUFF1_86 (N771, dN301);
buf BUFF1_87 (N774, dN297);
buf BUFF1_88 (N777, dN309);
buf BUFF1_89 (N780, dN305);
buf BUFF1_90 (N783, dN316);
buf BUFF1_91 (N786, dN313);
not NOT1_92 (dN792, N485);
not NOT1_93 (dN799, N495);
not NOT1_94 (N800, N499);
buf BUFF1_95 (dN805, N500);
nand NAND2_96 (N900, dN331, N606);
nand NAND2_97 (N901, dN328, N607);
nand NAND2_98 (N902, dN337, N608);
nand NAND2_99 (N903, dN334, N609);
nand NAND2_100 (N904, dN343, N610);
nand NAND2_101 (N905, dN340, N611);
nand NAND2_102 (N998, dN349, N733);
nand NAND2_103 (N999, dN346, N734);
and AND2_104 (dN1026, dN94, N500);
and AND2_105 (N1027, dN325, N651);
not NOT1_106 (dN1028, N651);
nand NAND2_107 (dN1029, dN231, N651);
not NOT1_108 (N1032, N544);
not NOT1_109 (N1033, N547);
and AND2_110 (N1034, N547, N544);
buf BUFF1_111 (N1037, N503);
not NOT1_112 (N1042, N509);
not NOT1_113 (N1053, N521);
and AND3_114 (N1064, dN80, N509, N521);
and AND3_115 (N1065, dN68, N509, N521);
and AND3_116 (N1066, dN79, N509, N521);
and AND3_117 (N1067, dN78, N509, N521);
and AND3_118 (N1068, dN77, N509, N521);
and AND2_119 (N1069, dN11, N537);
buf BUFF1_120 (N1070, N503);
not NOT1_121 (N1075, N550);
not NOT1_122 (N1086, N562);
and AND3_123 (N1097, dN76, N550, N562);
and AND3_124 (N1098, dN75, N550, N562);
and AND3_125 (N1099, dN74, N550, N562);
and AND3_126 (N1100, dN73, N550, N562);
and AND3_127 (N1101, dN72, N550, N562);
not NOT1_128 (N1102, N582);
not NOT1_129 (N1113, N594);
and AND3_130 (N1124, dN114, N582, N594);
and AND3_131 (N1125, dN113, N582, N594);
and AND3_132 (N1126, dN112, N582, N594);
and AND3_133 (N1127, dN111, N582, N594);
and AND2_134 (N1128, N582, N594);
nand NAND2_135 (N1129, N900, N901);
nand NAND2_136 (N1133, N902, N903);
nand NAND2_137 (N1137, N904, N905);
not NOT1_138 (N1140, N741);
nand NAND2_139 (N1141, N741, N612);
not NOT1_140 (N1142, N744);
not NOT1_141 (N1143, N747);
not NOT1_142 (N1144, N750);
not NOT1_143 (N1145, N753);
not NOT1_144 (N1146, N613);
not NOT1_145 (N1157, N625);
and AND3_146 (N1168, dN118, N613, N625);
and AND3_147 (N1169, dN107, N613, N625);
and AND3_148 (N1170, dN117, N613, N625);
and AND3_149 (N1171, dN116, N613, N625);
and AND3_150 (N1172, dN115, N613, N625);
not NOT1_151 (N1173, N637);
not NOT1_152 (N1178, N643);
not NOT1_153 (N1184, N768);
nand NAND2_154 (N1185, N768, N650);
not NOT1_155 (N1186, N771);
not NOT1_156 (N1187, N774);
not NOT1_157 (N1188, N777);
not NOT1_158 (N1189, N780);
buf BUFF1_159 (N1190, N506);
buf BUFF1_160 (N1195, N506);
not NOT1_161 (N1200, N693);
not NOT1_162 (N1205, N699);
not NOT1_163 (N1210, N735);
not NOT1_164 (N1211, N738);
not NOT1_165 (N1212, N756);
not NOT1_166 (N1213, N759);
not NOT1_167 (N1214, N762);
not NOT1_168 (N1215, N765);
nand NAND2_169 (N1216, N998, N999);
buf BUFF1_170 (N1219, N574);
buf BUFF1_171 (N1222, N578);
buf BUFF1_172 (N1225, N655);
buf BUFF1_173 (N1228, N659);
buf BUFF1_174 (N1231, N663);
buf BUFF1_175 (N1234, N667);
buf BUFF1_176 (N1237, N671);
buf BUFF1_177 (N1240, N675);
buf BUFF1_178 (N1243, N679);
buf BUFF1_179 (N1246, N683);
not NOT1_180 (N1249, N783);
not NOT1_181 (N1250, N786);
buf BUFF1_182 (N1251, N687);
buf BUFF1_183 (N1254, N705);
buf BUFF1_184 (N1257, N711);
buf BUFF1_185 (N1260, N715);
buf BUFF1_186 (N1263, N719);
buf BUFF1_187 (N1266, N723);
not NOT1_188 (dN1269, N1027);
and AND2_189 (N1275, dN325, N1032);
and AND2_190 (N1276, dN231, N1033);
buf BUFF1_191 (dN1277, N1034);
or OR2_192 (N1302, N1069, N543);
nand NAND2_193 (N1351, dN352, N1140);
nand NAND2_194 (N1352, N747, N1142);
nand NAND2_195 (N1353, N744, N1143);
nand NAND2_196 (N1354, N753, N1144);
nand NAND2_197 (N1355, N750, N1145);
nand NAND2_198 (N1395, dN355, N1184);
nand NAND2_199 (N1396, N774, N1186);
nand NAND2_200 (N1397, N771, N1187);
nand NAND2_201 (N1398, N780, N1188);
nand NAND2_202 (N1399, N777, N1189);
nand NAND2_203 (N1422, N738, N1210);
nand NAND2_204 (N1423, N735, N1211);
nand NAND2_205 (N1424, N759, N1212);
nand NAND2_206 (N1425, N756, N1213);
nand NAND2_207 (N1426, N765, N1214);
nand NAND2_208 (N1427, N762, N1215);
nand NAND2_209 (N1440, N786, N1249);
nand NAND2_210 (N1441, N783, N1250);
not NOT1_211 (dN1448, N1034);
not NOT1_212 (N1449, N1275);
not NOT1_213 (N1450, N1276);
and AND3_214 (N1451, dN93, N1042, N1053);
and AND3_215 (N1452, dN55, N509, N1053);
and AND3_216 (N1453, dN67, N1042, N521);
and AND3_217 (N1454, dN81, N1042, N1053);
and AND3_218 (N1455, dN43, N509, N1053);
and AND3_219 (N1456, dN56, N1042, N521);
and AND3_220 (N1457, dN92, N1042, N1053);
and AND3_221 (N1458, dN54, N509, N1053);
and AND3_222 (N1459, dN66, N1042, N521);
and AND3_223 (N1460, dN91, N1042, N1053);
and AND3_224 (N1461, dN53, N509, N1053);
and AND3_225 (N1462, dN65, N1042, N521);
and AND3_226 (N1463, dN90, N1042, N1053);
and AND3_227 (N1464, dN52, N509, N1053);
and AND3_228 (N1465, dN64, N1042, N521);
and AND3_229 (N1466, dN89, N1075, N1086);
and AND3_230 (N1467, dN51, N550, N1086);
and AND3_231 (N1468, dN63, N1075, N562);
and AND3_232 (N1469, dN88, N1075, N1086);
and AND3_233 (N1470, dN50, N550, N1086);
and AND3_234 (N1471, dN62, N1075, N562);
and AND3_235 (N1472, dN87, N1075, N1086);
and AND3_236 (N1473, dN49, N550, N1086);
and AND2_237 (N1474, N1075, N562);
and AND3_238 (N1475, dN86, N1075, N1086);
and AND3_239 (N1476, dN48, N550, N1086);
and AND3_240 (N1477, dN61, N1075, N562);
and AND3_241 (N1478, dN85, N1075, N1086);
and AND3_242 (N1479, dN47, N550, N1086);
and AND3_243 (N1480, dN60, N1075, N562);
and AND3_244 (N1481, dN138, N1102, N1113);
and AND3_245 (N1482, dN102, N582, N1113);
and AND3_246 (N1483, dN126, N1102, N594);
and AND3_247 (N1484, dN137, N1102, N1113);
and AND3_248 (N1485, dN101, N582, N1113);
and AND3_249 (N1486, dN125, N1102, N594);
and AND3_250 (N1487, dN136, N1102, N1113);
and AND3_251 (N1488, dN100, N582, N1113);
and AND3_252 (N1489, dN124, N1102, N594);
and AND3_253 (N1490, dN135, N1102, N1113);
and AND3_254 (N1491, dN99, N582, N1113);
and AND3_255 (N1492, dN123, N1102, N594);
and AND2_256 (N1493, N1102, N1113);
and AND2_257 (N1494, N582, N1113);
and AND2_258 (N1495, N1102, N594);
not NOT1_259 (N1496, N1129);
not NOT1_260 (N1499, N1133);
nand NAND2_261 (N1502, N1351, N1141);
nand NAND2_262 (N1506, N1352, N1353);
nand NAND2_263 (N1510, N1354, N1355);
buf BUFF1_264 (N1513, N1137);
buf BUFF1_265 (N1516, N1137);
not NOT1_266 (N1519, N1219);
not NOT1_267 (N1520, N1222);
not NOT1_268 (N1521, N1225);
not NOT1_269 (N1522, N1228);
not NOT1_270 (N1523, N1231);
not NOT1_271 (N1524, N1234);
not NOT1_272 (N1525, N1237);
not NOT1_273 (N1526, N1240);
not NOT1_274 (N1527, N1243);
not NOT1_275 (N1528, N1246);
and AND3_276 (N1529, dN142, N1146, N1157);
and AND3_277 (N1530, dN106, N613, N1157);
and AND3_278 (N1531, dN130, N1146, N625);
and AND3_279 (N1532, dN131, N1146, N1157);
and AND3_280 (N1533, dN95, N613, N1157);
and AND3_281 (N1534, dN119, N1146, N625);
and AND3_282 (N1535, dN141, N1146, N1157);
and AND3_283 (N1536, dN105, N613, N1157);
and AND3_284 (N1537, dN129, N1146, N625);
and AND3_285 (N1538, dN140, N1146, N1157);
and AND3_286 (N1539, dN104, N613, N1157);
and AND3_287 (N1540, dN128, N1146, N625);
and AND3_288 (N1541, dN139, N1146, N1157);
and AND3_289 (N1542, dN103, N613, N1157);
and AND3_290 (N1543, dN127, N1146, N625);
and AND2_291 (N1544, dN19, N1173);
and AND2_292 (N1545, dN4, N1173);
and AND2_293 (N1546, dN20, N1173);
and AND2_294 (N1547, dN5, N1173);
and AND2_295 (N1548, dN21, N1178);
and AND2_296 (N1549, dN22, N1178);
and AND2_297 (N1550, dN23, N1178);
and AND2_298 (N1551, dN6, N1178);
and AND2_299 (N1552, dN24, N1178);
nand NAND2_300 (N1553, N1395, N1185);
nand NAND2_301 (N1557, N1396, N1397);
nand NAND2_302 (N1561, N1398, N1399);
and AND2_303 (N1564, dN25, N1200);
and AND2_304 (N1565, dN32, N1200);
and AND2_305 (N1566, dN26, N1200);
and AND2_306 (N1567, dN33, N1200);
and AND2_307 (N1568, dN27, N1205);
and AND2_308 (N1569, dN34, N1205);
and AND2_309 (N1570, dN35, N1205);
and AND2_310 (N1571, dN28, N1205);
not NOT1_311 (N1572, N1251);
not NOT1_312 (N1573, N1254);
not NOT1_313 (N1574, N1257);
not NOT1_314 (N1575, N1260);
not NOT1_315 (N1576, N1263);
not NOT1_316 (N1577, N1266);
nand NAND2_317 (N1578, N1422, N1423);
not NOT1_318 (N1581, N1216);
nand NAND2_319 (N1582, N1426, N1427);
nand NAND2_320 (N1585, N1424, N1425);
nand NAND2_321 (N1588, N1440, N1441);
and AND2_322 (N1591, N1449, N1450);
or OR4_323 (N1596, N1451, N1452, N1453, N1064);
or OR4_324 (N1600, N1454, N1455, N1456, N1065);
or OR4_325 (N1606, N1457, N1458, N1459, N1066);
or OR4_326 (N1612, N1460, N1461, N1462, N1067);
or OR4_327 (N1615, N1463, N1464, N1465, N1068);
or OR4_328 (N1619, N1466, N1467, N1468, N1097);
or OR4_329 (N1624, N1469, N1470, N1471, N1098);
or OR4_330 (N1628, N1472, N1473, N1474, N1099);
or OR4_331 (N1631, N1475, N1476, N1477, N1100);
or OR4_332 (N1634, N1478, N1479, N1480, N1101);
or OR4_333 (N1637, N1481, N1482, N1483, N1124);
or OR4_334 (N1642, N1484, N1485, N1486, N1125);
or OR4_335 (N1647, N1487, N1488, N1489, N1126);
or OR4_336 (N1651, N1490, N1491, N1492, N1127);
or OR4_337 (N1656, N1493, N1494, N1495, N1128);
or OR4_338 (N1676, N1532, N1533, N1534, N1169);
or OR4_339 (N1681, N1535, N1536, N1537, N1170);
or OR4_340 (N1686, N1538, N1539, N1540, N1171);
or OR4_341 (N1690, N1541, N1542, N1543, N1172);
or OR4_342 (N1708, N1529, N1530, N1531, N1168);
buf BUFF1_343 (dN1726, N1591);
not NOT1_344 (N1770, N1502);
not NOT1_345 (N1773, N1506);
not NOT1_346 (N1776, N1513);
not NOT1_347 (N1777, N1516);
buf BUFF1_348 (N1778, N1510);
buf BUFF1_349 (N1781, N1510);
and AND3_350 (N1784, N1133, N1129, N1513);
and AND3_351 (N1785, N1499, N1496, N1516);
not NOT1_352 (N1795, N1553);
not NOT1_353 (N1798, N1557);
buf BUFF1_354 (N1801, N1561);
buf BUFF1_355 (N1804, N1561);
not NOT1_356 (N1807, N1588);
not NOT1_357 (N1808, N1578);
nand NAND2_358 (N1809, N1578, N1581);
not NOT1_359 (N1810, N1582);
not NOT1_360 (N1811, N1585);
and AND2_361 (N1813, N1596, dN241);
and AND2_362 (N1814, N1606, dN241);
and AND2_363 (N1815, N1600, dN241);
not NOT1_364 (dN1816, N1642);
not NOT1_365 (dN1817, N1647);
not NOT1_366 (dN1818, N1637);
not NOT1_367 (dN1819, N1624);
not NOT1_368 (dN1820, N1619);
not NOT1_369 (dN1821, N1615);
and AND4_370 (N1822, N496, dN224, dN36, N1591);
and AND4_371 (N1823, N496, dN224, N1591, N486);
buf BUFF1_372 (N1824, N1596);
not NOT1_373 (N1827, N1606);
and AND2_374 (N1830, N1600, N537);
and AND2_375 (N1831, N1606, N537);
and AND2_376 (N1832, N1619, dN246);
not NOT1_377 (N1833, N1596);
not NOT1_378 (N1836, N1600);
not NOT1_379 (N1841, N1606);
buf BUFF1_380 (N1848, N1612);
buf BUFF1_381 (N1852, N1615);
buf BUFF1_382 (N1856, N1619);
buf BUFF1_383 (N1863, N1624);
buf BUFF1_384 (N1870, N1628);
buf BUFF1_385 (N1875, N1631);
buf BUFF1_386 (N1880, N1634);
nand NAND2_387 (N1885, N727, N1651);
nand NAND2_388 (N1888, N730, N1656);
buf BUFF1_389 (N1891, N1686);
and AND2_390 (N1894, N1637, N425);
not NOT1_391 (N1897, N1642);
and AND3_392 (N1908, N1496, N1133, N1776);
and AND3_393 (N1909, N1129, N1499, N1777);
and AND2_394 (N1910, N1600, N637);
and AND2_395 (N1911, N1606, N637);
and AND2_396 (N1912, N1612, N637);
and AND2_397 (N1913, N1615, N637);
and AND2_398 (N1914, N1619, N643);
and AND2_399 (N1915, N1624, N643);
and AND2_400 (N1916, N1628, N643);
and AND2_401 (N1917, N1631, N643);
and AND2_402 (N1918, N1634, N643);
not NOT1_403 (N1919, N1708);
and AND2_404 (N1928, N1676, N693);
and AND2_405 (N1929, N1681, N693);
and AND2_406 (N1930, N1686, N693);
and AND2_407 (N1931, N1690, N693);
and AND2_408 (N1932, N1637, N699);
and AND2_409 (N1933, N1642, N699);
and AND2_410 (N1934, N1647, N699);
and AND2_411 (N1935, N1651, N699);
buf BUFF1_412 (N1936, N1600);
nand NAND2_413 (N1939, N1216, N1808);
nand NAND2_414 (N1940, N1585, N1810);
nand NAND2_415 (N1941, N1582, N1811);
buf BUFF1_416 (N1942, N1676);
buf BUFF1_417 (N1945, N1686);
buf BUFF1_418 (N1948, N1681);
buf BUFF1_419 (N1951, N1637);
buf BUFF1_420 (N1954, N1690);
buf BUFF1_421 (N1957, N1647);
buf BUFF1_422 (N1960, N1642);
buf BUFF1_423 (N1963, N1656);
buf BUFF1_424 (N1966, N1651);
or OR2_425 (dN1969, N533, N1815);
not NOT1_426 (dN1970, N1822);
not NOT1_427 (dN1971, N1823);
buf BUFF1_428 (dN2010, N1848);
buf BUFF1_429 (dN2012, N1852);
buf BUFF1_430 (dN2014, N1856);
buf BUFF1_431 (dN2016, N1863);
buf BUFF1_432 (dN2018, N1870);
buf BUFF1_433 (dN2020, N1875);
buf BUFF1_434 (dN2022, N1880);
not NOT1_435 (N2028, N1778);
not NOT1_436 (N2029, N1781);
nor NOR2_437 (N2030, N1908, N1784);
nor NOR2_438 (N2031, N1909, N1785);
and AND3_439 (N2032, N1506, N1502, N1778);
and AND3_440 (N2033, N1773, N1770, N1781);
or OR2_441 (N2034, N1571, N1935);
not NOT1_442 (N2040, N1801);
not NOT1_443 (N2041, N1804);
and AND3_444 (N2042, N1557, N1553, N1801);
and AND3_445 (N2043, N1798, N1795, N1804);
nand NAND2_446 (N2046, N1939, N1809);
nand NAND2_447 (N2049, N1940, N1941);
or OR2_448 (N2052, N1544, N1910);
or OR2_449 (N2055, N1545, N1911);
or OR2_450 (N2058, N1546, N1912);
or OR2_451 (N2061, N1547, N1913);
or OR2_452 (N2064, N1548, N1914);
or OR2_453 (N2067, N1549, N1915);
or OR2_454 (N2070, N1550, N1916);
or OR2_455 (N2073, N1551, N1917);
or OR2_456 (N2076, N1552, N1918);
or OR2_457 (N2079, N1564, N1928);
or OR2_458 (N2095, N1565, N1929);
or OR2_459 (N2098, N1566, N1930);
or OR2_460 (N2101, N1567, N1931);
or OR2_461 (N2104, N1568, N1932);
or OR2_462 (N2107, N1569, N1933);
or OR2_463 (N2110, N1570, N1934);
and AND3_464 (N2113, N1897, N1894, dN40);
not NOT1_465 (N2119, N1894);
nand NAND2_466 (N2120, N408, N1827);
and AND2_467 (N2125, N1824, N537);
and AND2_468 (N2126, N1852, dN246);
and AND2_469 (N2127, N1848, N537);
not NOT1_470 (N2128, N1848);
not NOT1_471 (N2135, N1852);
not NOT1_472 (N2141, N1863);
not NOT1_473 (N2144, N1870);
not NOT1_474 (N2147, N1875);
not NOT1_475 (N2150, N1880);
and AND2_476 (N2153, N727, N1885);
and AND2_477 (N2154, N1885, N1651);
and AND2_478 (N2155, N730, N1888);
and AND2_479 (N2156, N1888, N1656);
and AND3_480 (N2157, N1770, N1506, N2028);
and AND3_481 (N2158, N1502, N1773, N2029);
not NOT1_482 (N2171, N1942);
nand NAND2_483 (N2172, N1942, N1919);
not NOT1_484 (N2173, N1945);
not NOT1_485 (N2174, N1948);
not NOT1_486 (N2175, N1951);
not NOT1_487 (N2176, N1954);
and AND3_488 (N2177, N1795, N1557, N2040);
and AND3_489 (N2178, N1553, N1798, N2041);
buf BUFF1_490 (N2185, N1836);
buf BUFF1_491 (N2188, N1833);
buf BUFF1_492 (N2191, N1841);
not NOT1_493 (N2194, N1856);
not NOT1_494 (N2197, N1827);
not NOT1_495 (N2200, N1936);
buf BUFF1_496 (N2201, N1836);
buf BUFF1_497 (N2204, N1833);
buf BUFF1_498 (N2207, N1841);
buf BUFF1_499 (N2210, N1824);
buf BUFF1_500 (N2213, N1841);
buf BUFF1_501 (N2216, N1841);
nand NAND2_502 (N2219, N2031, N2030);
not NOT1_503 (N2234, N1957);
not NOT1_504 (N2235, N1960);
not NOT1_505 (N2236, N1963);
not NOT1_506 (N2237, N1966);
and AND3_507 (N2250, dN40, N1897, N2119);
or OR2_508 (N2266, N1831, N2126);
or OR2_509 (N2269, N2127, N1832);
or OR2_510 (N2291, N2153, N2154);
or OR2_511 (N2294, N2155, N2156);
nor NOR2_512 (N2297, N2157, N2032);
nor NOR2_513 (N2298, N2158, N2033);
not NOT1_514 (N2300, N2046);
not NOT1_515 (N2301, N2049);
nand NAND2_516 (N2302, N2052, N1519);
not NOT1_517 (N2303, N2052);
nand NAND2_518 (N2304, N2055, N1520);
not NOT1_519 (N2305, N2055);
nand NAND2_520 (N2306, N2058, N1521);
not NOT1_521 (N2307, N2058);
nand NAND2_522 (N2308, N2061, N1522);
not NOT1_523 (N2309, N2061);
nand NAND2_524 (N2310, N2064, N1523);
not NOT1_525 (N2311, N2064);
nand NAND2_526 (N2312, N2067, N1524);
not NOT1_527 (N2313, N2067);
nand NAND2_528 (N2314, N2070, N1525);
not NOT1_529 (N2315, N2070);
nand NAND2_530 (N2316, N2073, N1526);
not NOT1_531 (N2317, N2073);
nand NAND2_532 (N2318, N2076, N1527);
not NOT1_533 (N2319, N2076);
nand NAND2_534 (N2320, N2079, N1528);
not NOT1_535 (N2321, N2079);
nand NAND2_536 (N2322, N1708, N2171);
nand NAND2_537 (N2323, N1948, N2173);
nand NAND2_538 (N2324, N1945, N2174);
nand NAND2_539 (N2325, N1954, N2175);
nand NAND2_540 (N2326, N1951, N2176);
nor NOR2_541 (N2327, N2177, N2042);
nor NOR2_542 (N2328, N2178, N2043);
nand NAND2_543 (N2329, N2095, N1572);
not NOT1_544 (N2330, N2095);
nand NAND2_545 (N2331, N2098, N1573);
not NOT1_546 (N2332, N2098);
nand NAND2_547 (N2333, N2101, N1574);
not NOT1_548 (N2334, N2101);
nand NAND2_549 (N2335, N2104, N1575);
not NOT1_550 (N2336, N2104);
nand NAND2_551 (N2337, N2107, N1576);
not NOT1_552 (N2338, N2107);
nand NAND2_553 (N2339, N2110, N1577);
not NOT1_554 (N2340, N2110);
nand NAND2_555 (N2354, N1960, N2234);
nand NAND2_556 (N2355, N1957, N2235);
nand NAND2_557 (N2356, N1966, N2236);
nand NAND2_558 (N2357, N1963, N2237);
and AND2_559 (N2358, N2120, N533);
not NOT1_560 (N2359, N2113);
not NOT1_561 (N2364, N2185);
not NOT1_562 (N2365, N2188);
not NOT1_563 (N2366, N2191);
not NOT1_564 (N2367, N2194);
buf BUFF1_565 (N2368, N2120);
not NOT1_566 (N2372, N2201);
not NOT1_567 (N2373, N2204);
not NOT1_568 (N2374, N2207);
not NOT1_569 (N2375, N2210);
not NOT1_570 (N2376, N2213);
not NOT1_571 (N2377, N2113);
buf BUFF1_572 (N2382, N2113);
and AND2_573 (N2386, N2120, dN246);
buf BUFF1_574 (dN2387, N2266);
buf BUFF1_575 (dN2388, N2266);
buf BUFF1_576 (dN2389, N2269);
buf BUFF1_577 (dN2390, N2269);
buf BUFF1_578 (N2391, N2113);
not NOT1_579 (N2395, N2113);
nand NAND2_580 (N2400, N2219, N2300);
not NOT1_581 (N2403, N2216);
not NOT1_582 (N2406, N2219);
nand NAND2_583 (N2407, N1219, N2303);
nand NAND2_584 (N2408, N1222, N2305);
nand NAND2_585 (N2409, N1225, N2307);
nand NAND2_586 (N2410, N1228, N2309);
nand NAND2_587 (N2411, N1231, N2311);
nand NAND2_588 (N2412, N1234, N2313);
nand NAND2_589 (N2413, N1237, N2315);
nand NAND2_590 (N2414, N1240, N2317);
nand NAND2_591 (N2415, N1243, N2319);
nand NAND2_592 (N2416, N1246, N2321);
nand NAND2_593 (N2417, N2322, N2172);
nand NAND2_594 (N2421, N2323, N2324);
nand NAND2_595 (N2425, N2325, N2326);
nand NAND2_596 (N2428, N1251, N2330);
nand NAND2_597 (N2429, N1254, N2332);
nand NAND2_598 (N2430, N1257, N2334);
nand NAND2_599 (N2431, N1260, N2336);
nand NAND2_600 (N2432, N1263, N2338);
nand NAND2_601 (N2433, N1266, N2340);
buf BUFF1_602 (N2434, N2128);
buf BUFF1_603 (N2437, N2135);
buf BUFF1_604 (N2440, N2144);
buf BUFF1_605 (N2443, N2141);
buf BUFF1_606 (N2446, N2150);
buf BUFF1_607 (N2449, N2147);
not NOT1_608 (N2452, N2197);
nand NAND2_609 (N2453, N2197, N2200);
buf BUFF1_610 (N2454, N2128);
buf BUFF1_611 (N2457, N2144);
buf BUFF1_612 (N2460, N2141);
buf BUFF1_613 (N2463, N2150);
buf BUFF1_614 (N2466, N2147);
not NOT1_615 (N2469, N2120);
buf BUFF1_616 (N2472, N2128);
buf BUFF1_617 (N2475, N2135);
buf BUFF1_618 (N2478, N2128);
buf BUFF1_619 (N2481, N2135);
nand NAND2_620 (N2484, N2298, N2297);
nand NAND2_621 (N2487, N2356, N2357);
nand NAND2_622 (N2490, N2354, N2355);
nand NAND2_623 (N2493, N2328, N2327);
or OR2_624 (dN2496, N2358, N1814);
nand NAND2_625 (N2503, N2188, N2364);
nand NAND2_626 (N2504, N2185, N2365);
nand NAND2_627 (N2510, N2204, N2372);
nand NAND2_628 (N2511, N2201, N2373);
or OR2_629 (N2521, N1830, N2386);
nand NAND2_630 (N2528, N2046, N2406);
not NOT1_631 (N2531, N2291);
not NOT1_632 (N2534, N2294);
buf BUFF1_633 (N2537, N2250);
buf BUFF1_634 (N2540, N2250);
nand NAND2_635 (N2544, N2302, N2407);
nand NAND2_636 (N2545, N2304, N2408);
nand NAND2_637 (N2546, N2306, N2409);
nand NAND2_638 (N2547, N2308, N2410);
nand NAND2_639 (N2548, N2310, N2411);
nand NAND2_640 (N2549, N2312, N2412);
nand NAND2_641 (N2550, N2314, N2413);
nand NAND2_642 (N2551, N2316, N2414);
nand NAND2_643 (N2552, N2318, N2415);
nand NAND2_644 (N2553, N2320, N2416);
nand NAND2_645 (N2563, N2329, N2428);
nand NAND2_646 (N2564, N2331, N2429);
nand NAND2_647 (N2565, N2333, N2430);
nand NAND2_648 (N2566, N2335, N2431);
nand NAND2_649 (N2567, N2337, N2432);
nand NAND2_650 (N2568, N2339, N2433);
nand NAND2_651 (N2579, N1936, N2452);
buf BUFF1_652 (N2603, N2359);
and AND2_653 (N2607, N1880, N2377);
and AND2_654 (N2608, N1676, N2377);
and AND2_655 (N2609, N1681, N2377);
and AND2_656 (N2610, N1891, N2377);
and AND2_657 (N2611, N1856, N2382);
and AND2_658 (N2612, N1863, N2382);
nand NAND2_659 (N2613, N2503, N2504);
not NOT1_660 (N2617, N2434);
nand NAND2_661 (N2618, N2434, N2366);
nand NAND2_662 (N2619, N2437, N2367);
not NOT1_663 (N2620, N2437);
not NOT1_664 (N2621, N2368);
nand NAND2_665 (N2624, N2510, N2511);
not NOT1_666 (N2628, N2454);
nand NAND2_667 (N2629, N2454, N2374);
not NOT1_668 (N2630, N2472);
and AND2_669 (N2631, N1856, N2391);
and AND2_670 (N2632, N1863, N2391);
and AND2_671 (N2633, N1880, N2395);
and AND2_672 (N2634, N1676, N2395);
and AND2_673 (N2635, N1681, N2395);
and AND2_674 (N2636, N1891, N2395);
not NOT1_675 (N2638, N2382);
buf BUFF1_676 (dN2643, N2521);
buf BUFF1_677 (dN2644, N2521);
not NOT1_678 (N2645, N2475);
not NOT1_679 (N2646, N2391);
nand NAND2_680 (N2652, N2528, N2400);
not NOT1_681 (N2655, N2478);
not NOT1_682 (N2656, N2481);
buf BUFF1_683 (N2659, N2359);
not NOT1_684 (N2663, N2484);
nand NAND2_685 (N2664, N2484, N2301);
not NOT1_686 (N2665, N2553);
not NOT1_687 (N2666, N2552);
not NOT1_688 (N2667, N2551);
not NOT1_689 (N2668, N2550);
not NOT1_690 (N2669, N2549);
not NOT1_691 (N2670, N2548);
not NOT1_692 (N2671, N2547);
not NOT1_693 (N2672, N2546);
not NOT1_694 (N2673, N2545);
not NOT1_695 (N2674, N2544);
not NOT1_696 (N2675, N2568);
not NOT1_697 (N2676, N2567);
not NOT1_698 (N2677, N2566);
not NOT1_699 (N2678, N2565);
not NOT1_700 (N2679, N2564);
not NOT1_701 (N2680, N2563);
not NOT1_702 (N2681, N2417);
not NOT1_703 (N2684, N2421);
buf BUFF1_704 (N2687, N2425);
buf BUFF1_705 (N2690, N2425);
not NOT1_706 (N2693, N2493);
nand NAND2_707 (N2694, N2493, N1807);
not NOT1_708 (N2695, N2440);
not NOT1_709 (N2696, N2443);
not NOT1_710 (N2697, N2446);
not NOT1_711 (N2698, N2449);
not NOT1_712 (N2699, N2457);
not NOT1_713 (N2700, N2460);
not NOT1_714 (N2701, N2463);
not NOT1_715 (N2702, N2466);
nand NAND2_716 (N2703, N2579, N2453);
not NOT1_717 (N2706, N2469);
not NOT1_718 (N2707, N2487);
not NOT1_719 (N2708, N2490);
and AND2_720 (N2709, N2294, N2534);
and AND2_721 (N2710, N2291, N2531);
nand NAND2_722 (N2719, N2191, N2617);
nand NAND2_723 (N2720, N2194, N2620);
nand NAND2_724 (N2726, N2207, N2628);
buf BUFF1_725 (N2729, N2537);
buf BUFF1_726 (N2738, N2537);
not NOT1_727 (N2743, N2652);
nand NAND2_728 (N2747, N2049, N2663);
and AND5_729 (N2748, N2665, N2666, N2667, N2668, N2669);
and AND5_730 (N2749, N2670, N2671, N2672, N2673, N2674);
and AND2_731 (N2750, N2034, N2675);
and AND5_732 (N2751, N2676, N2677, N2678, N2679, N2680);
nand NAND2_733 (N2760, N1588, N2693);
buf BUFF1_734 (N2761, N2540);
buf BUFF1_735 (N2766, N2540);
nand NAND2_736 (N2771, N2443, N2695);
nand NAND2_737 (N2772, N2440, N2696);
nand NAND2_738 (N2773, N2449, N2697);
nand NAND2_739 (N2774, N2446, N2698);
nand NAND2_740 (N2775, N2460, N2699);
nand NAND2_741 (N2776, N2457, N2700);
nand NAND2_742 (N2777, N2466, N2701);
nand NAND2_743 (N2778, N2463, N2702);
nand NAND2_744 (N2781, N2490, N2707);
nand NAND2_745 (N2782, N2487, N2708);
or OR2_746 (N2783, N2709, N2534);
or OR2_747 (N2784, N2710, N2531);
and AND2_748 (N2789, N1856, N2638);
and AND2_749 (N2790, N1863, N2638);
and AND2_750 (N2791, N1870, N2638);
and AND2_751 (N2792, N1875, N2638);
not NOT1_752 (N2793, N2613);
nand NAND2_753 (N2796, N2719, N2618);
nand NAND2_754 (N2800, N2619, N2720);
not NOT1_755 (N2803, N2624);
nand NAND2_756 (N2806, N2726, N2629);
and AND2_757 (N2809, N1856, N2646);
and AND2_758 (N2810, N1863, N2646);
and AND2_759 (N2811, N1870, N2646);
and AND2_760 (N2812, N1875, N2646);
and AND2_761 (N2817, N2743, dN14);
buf BUFF1_762 (N2820, N2603);
nand NAND2_763 (N2826, N2747, N2664);
and AND2_764 (N2829, N2748, N2749);
and AND2_765 (N2830, N2750, N2751);
buf BUFF1_766 (N2831, N2659);
not NOT1_767 (N2837, N2687);
not NOT1_768 (N2838, N2690);
and AND3_769 (N2839, N2421, N2417, N2687);
and AND3_770 (N2840, N2684, N2681, N2690);
nand NAND2_771 (N2841, N2760, N2694);
buf BUFF1_772 (N2844, N2603);
buf BUFF1_773 (N2854, N2603);
buf BUFF1_774 (N2859, N2659);
buf BUFF1_775 (N2869, N2659);
nand NAND2_776 (N2874, N2773, N2774);
nand NAND2_777 (N2877, N2771, N2772);
not NOT1_778 (N2880, N2703);
nand NAND2_779 (N2881, N2703, N2706);
nand NAND2_780 (N2882, N2777, N2778);
nand NAND2_781 (N2885, N2775, N2776);
nand NAND2_782 (N2888, N2781, N2782);
nand NAND2_783 (dN2891, N2783, N2784);
and AND2_784 (N2894, N2607, N2729);
and AND2_785 (N2895, N2608, N2729);
and AND2_786 (N2896, N2609, N2729);
and AND2_787 (N2897, N2610, N2729);
or OR2_788 (N2898, N2789, N2611);
or OR2_789 (N2899, N2790, N2612);
and AND2_790 (N2900, N2791, N1037);
and AND2_791 (N2901, N2792, N1037);
or OR2_792 (N2914, N2809, N2631);
or OR2_793 (N2915, N2810, N2632);
and AND2_794 (N2916, N2811, N1070);
and AND2_795 (N2917, N2812, N1070);
and AND2_796 (N2918, N2633, N2738);
and AND2_797 (N2919, N2634, N2738);
and AND2_798 (N2920, N2635, N2738);
and AND2_799 (N2921, N2636, N2738);
buf BUFF1_800 (dN2925, N2817);
and AND3_801 (N2931, N2829, N2830, N1302);
and AND3_802 (N2938, N2681, N2421, N2837);
and AND3_803 (N2939, N2417, N2684, N2838);
nand NAND2_804 (N2963, N2469, N2880);
not NOT1_805 (dN2970, N2841);
not NOT1_806 (dN2971, N2826);
not NOT1_807 (N2972, N2894);
not NOT1_808 (N2975, N2895);
not NOT1_809 (N2978, N2896);
not NOT1_810 (N2981, N2897);
and AND2_811 (N2984, N2898, N1037);
and AND2_812 (N2985, N2899, N1037);
not NOT1_813 (N2986, N2900);
not NOT1_814 (N2989, N2901);
not NOT1_815 (N2992, N2796);
buf BUFF1_816 (N2995, N2800);
buf BUFF1_817 (N2998, N2800);
buf BUFF1_818 (N3001, N2806);
buf BUFF1_819 (N3004, N2806);
and AND2_820 (N3007, N574, N2820);
and AND2_821 (N3008, N2914, N1070);
and AND2_822 (N3009, N2915, N1070);
not NOT1_823 (N3010, N2916);
not NOT1_824 (N3013, N2917);
not NOT1_825 (N3016, N2918);
not NOT1_826 (N3019, N2919);
not NOT1_827 (N3022, N2920);
not NOT1_828 (N3025, N2921);
not NOT1_829 (N3028, N2817);
and AND2_830 (N3029, N574, N2831);
not NOT1_831 (N3030, N2820);
and AND2_832 (N3035, N578, N2820);
and AND2_833 (N3036, N655, N2820);
and AND2_834 (N3037, N659, N2820);
buf BUFF1_835 (dN3038, N2931);
not NOT1_836 (N3039, N2831);
and AND2_837 (N3044, N578, N2831);
and AND2_838 (N3045, N655, N2831);
and AND2_839 (N3046, N659, N2831);
nor NOR2_840 (N3047, N2938, N2839);
nor NOR2_841 (N3048, N2939, N2840);
not NOT1_842 (N3049, N2888);
not NOT1_843 (N3050, N2844);
and AND2_844 (N3053, N663, N2844);
and AND2_845 (N3054, N667, N2844);
and AND2_846 (N3055, N671, N2844);
and AND2_847 (N3056, N675, N2844);
and AND2_848 (N3057, N679, N2854);
and AND2_849 (N3058, N683, N2854);
and AND2_850 (N3059, N687, N2854);
and AND2_851 (N3060, N705, N2854);
not NOT1_852 (N3061, N2859);
and AND2_853 (N3064, N663, N2859);
and AND2_854 (N3065, N667, N2859);
and AND2_855 (N3066, N671, N2859);
and AND2_856 (N3067, N675, N2859);
and AND2_857 (N3068, N679, N2869);
and AND2_858 (N3069, N683, N2869);
and AND2_859 (N3070, N687, N2869);
and AND2_860 (N3071, N705, N2869);
not NOT1_861 (N3072, N2874);
not NOT1_862 (N3073, N2877);
not NOT1_863 (N3074, N2882);
not NOT1_864 (N3075, N2885);
nand NAND2_865 (N3076, N2881, N2963);
not NOT1_866 (dN3079, N2931);
not NOT1_867 (N3088, N2984);
not NOT1_868 (N3091, N2985);
not NOT1_869 (N3110, N3008);
not NOT1_870 (N3113, N3009);
and AND2_871 (N3137, N3055, N1190);
and AND2_872 (N3140, N3056, N1190);
and AND2_873 (N3143, N3057, N2761);
and AND2_874 (N3146, N3058, N2761);
and AND2_875 (N3149, N3059, N2761);
and AND2_876 (N3152, N3060, N2761);
and AND2_877 (N3157, N3066, N1195);
and AND2_878 (N3160, N3067, N1195);
and AND2_879 (N3163, N3068, N2766);
and AND2_880 (N3166, N3069, N2766);
and AND2_881 (N3169, N3070, N2766);
and AND2_882 (N3172, N3071, N2766);
nand NAND2_883 (N3175, N2877, N3072);
nand NAND2_884 (N3176, N2874, N3073);
nand NAND2_885 (N3177, N2885, N3074);
nand NAND2_886 (N3178, N2882, N3075);
nand NAND2_887 (N3180, N3048, N3047);
not NOT1_888 (N3187, N2995);
not NOT1_889 (N3188, N2998);
not NOT1_890 (N3189, N3001);
not NOT1_891 (N3190, N3004);
and AND3_892 (N3191, N2796, N2613, N2995);
and AND3_893 (N3192, N2992, N2793, N2998);
and AND3_894 (N3193, N2624, N2368, N3001);
and AND3_895 (N3194, N2803, N2621, N3004);
nand NAND2_896 (N3195, N3076, N2375);
not NOT1_897 (N3196, N3076);
and AND2_898 (N3197, N687, N3030);
and AND2_899 (N3208, N687, N3039);
and AND2_900 (N3215, N705, N3030);
and AND2_901 (N3216, N711, N3030);
and AND2_902 (N3217, N715, N3030);
and AND2_903 (N3218, N705, N3039);
and AND2_904 (N3219, N711, N3039);
and AND2_905 (N3220, N715, N3039);
and AND2_906 (N3222, N719, N3050);
and AND2_907 (N3223, N723, N3050);
and AND2_908 (N3230, N719, N3061);
and AND2_909 (N3231, N723, N3061);
nand NAND2_910 (N3238, N3175, N3176);
nand NAND2_911 (N3241, N3177, N3178);
buf BUFF1_912 (N3244, N2981);
buf BUFF1_913 (N3247, N2978);
buf BUFF1_914 (N3250, N2975);
buf BUFF1_915 (N3253, N2972);
buf BUFF1_916 (N3256, N2989);
buf BUFF1_917 (N3259, N2986);
buf BUFF1_918 (N3262, N3025);
buf BUFF1_919 (N3265, N3022);
buf BUFF1_920 (N3268, N3019);
buf BUFF1_921 (N3271, N3016);
buf BUFF1_922 (N3274, N3013);
buf BUFF1_923 (N3277, N3010);
and AND3_924 (N3281, N2793, N2796, N3187);
and AND3_925 (N3282, N2613, N2992, N3188);
and AND3_926 (N3283, N2621, N2624, N3189);
and AND3_927 (N3284, N2368, N2803, N3190);
nand NAND2_928 (N3286, N2210, N3196);
or OR2_929 (N3288, N3197, N3007);
nand NAND2_930 (N3289, N3180, N3049);
and AND2_931 (N3291, N3152, N2981);
and AND2_932 (N3293, N3149, N2978);
and AND2_933 (N3295, N3146, N2975);
and AND2_934 (N3296, N2972, N3143);
and AND2_935 (N3299, N3140, N2989);
and AND2_936 (N3301, N3137, N2986);
or OR2_937 (N3302, N3208, N3029);
and AND2_938 (N3304, N3172, N3025);
and AND2_939 (N3306, N3169, N3022);
and AND2_940 (N3308, N3166, N3019);
and AND2_941 (N3309, N3016, N3163);
and AND2_942 (N3312, N3160, N3013);
and AND2_943 (N3314, N3157, N3010);
or OR2_944 (N3315, N3215, N3035);
or OR2_945 (N3318, N3216, N3036);
or OR2_946 (N3321, N3217, N3037);
or OR2_947 (N3324, N3218, N3044);
or OR2_948 (N3327, N3219, N3045);
or OR2_949 (N3330, N3220, N3046);
not NOT1_950 (N3333, N3180);
or OR2_951 (N3334, N3222, N3053);
or OR2_952 (N3335, N3223, N3054);
or OR2_953 (N3336, N3230, N3064);
or OR2_954 (N3337, N3231, N3065);
buf BUFF1_955 (N3340, N3152);
buf BUFF1_956 (N3344, N3149);
buf BUFF1_957 (N3348, N3146);
buf BUFF1_958 (N3352, N3143);
buf BUFF1_959 (N3356, N3140);
buf BUFF1_960 (N3360, N3137);
buf BUFF1_961 (N3364, N3091);
buf BUFF1_962 (N3367, N3088);
buf BUFF1_963 (N3370, N3172);
buf BUFF1_964 (N3374, N3169);
buf BUFF1_965 (N3378, N3166);
buf BUFF1_966 (N3382, N3163);
buf BUFF1_967 (N3386, N3160);
buf BUFF1_968 (N3390, N3157);
buf BUFF1_969 (N3394, N3113);
buf BUFF1_970 (N3397, N3110);
nand NAND2_971 (N3400, N3195, N3286);
nor NOR2_972 (N3401, N3281, N3191);
nor NOR2_973 (N3402, N3282, N3192);
nor NOR2_974 (N3403, N3283, N3193);
nor NOR2_975 (N3404, N3284, N3194);
not NOT1_976 (N3405, N3238);
not NOT1_977 (N3406, N3241);
and AND2_978 (N3409, N3288, N1836);
nand NAND2_979 (N3410, N2888, N3333);
not NOT1_980 (N3412, N3244);
not NOT1_981 (N3414, N3247);
not NOT1_982 (N3416, N3250);
not NOT1_983 (N3418, N3253);
not NOT1_984 (N3420, N3256);
not NOT1_985 (N3422, N3259);
and AND2_986 (N3428, N3302, N1836);
not NOT1_987 (N3430, N3262);
not NOT1_988 (N3432, N3265);
not NOT1_989 (N3434, N3268);
not NOT1_990 (N3436, N3271);
not NOT1_991 (N3438, N3274);
not NOT1_992 (N3440, N3277);
and AND2_993 (N3450, N3334, N1190);
and AND2_994 (N3453, N3335, N1190);
and AND2_995 (N3456, N3336, N1195);
and AND2_996 (N3459, N3337, N1195);
and AND2_997 (N3478, N3400, N533);
and AND2_998 (N3479, N3318, N2128);
and AND2_999 (N3480, N3315, N1841);
nand NAND2_1000 (N3481, N3410, N3289);
not NOT1_1001 (N3482, N3340);
nand NAND2_1002 (N3483, N3340, N3412);
not NOT1_1003 (N3484, N3344);
nand NAND2_1004 (N3485, N3344, N3414);
not NOT1_1005 (N3486, N3348);
nand NAND2_1006 (N3487, N3348, N3416);
not NOT1_1007 (N3488, N3352);
nand NAND2_1008 (N3489, N3352, N3418);
not NOT1_1009 (N3490, N3356);
nand NAND2_1010 (N3491, N3356, N3420);
not NOT1_1011 (N3492, N3360);
nand NAND2_1012 (N3493, N3360, N3422);
not NOT1_1013 (N3494, N3364);
not NOT1_1014 (N3496, N3367);
and AND2_1015 (N3498, N3321, N2135);
and AND2_1016 (N3499, N3327, N2128);
and AND2_1017 (N3500, N3324, N1841);
not NOT1_1018 (N3501, N3370);
nand NAND2_1019 (N3502, N3370, N3430);
not NOT1_1020 (N3503, N3374);
nand NAND2_1021 (N3504, N3374, N3432);
not NOT1_1022 (N3505, N3378);
nand NAND2_1023 (N3506, N3378, N3434);
not NOT1_1024 (N3507, N3382);
nand NAND2_1025 (N3508, N3382, N3436);
not NOT1_1026 (N3509, N3386);
nand NAND2_1027 (N3510, N3386, N3438);
not NOT1_1028 (N3511, N3390);
nand NAND2_1029 (N3512, N3390, N3440);
not NOT1_1030 (N3513, N3394);
not NOT1_1031 (N3515, N3397);
and AND2_1032 (N3517, N3330, N2135);
nand NAND2_1033 (N3522, N3402, N3401);
nand NAND2_1034 (N3525, N3404, N3403);
buf BUFF1_1035 (N3528, N3318);
buf BUFF1_1036 (N3531, N3315);
buf BUFF1_1037 (N3534, N3321);
buf BUFF1_1038 (N3537, N3327);
buf BUFF1_1039 (N3540, N3324);
buf BUFF1_1040 (N3543, N3330);
or OR2_1041 (dN3546, N3478, N1813);
not NOT1_1042 (N3551, N3481);
nand NAND2_1043 (N3552, N3244, N3482);
nand NAND2_1044 (N3553, N3247, N3484);
nand NAND2_1045 (N3554, N3250, N3486);
nand NAND2_1046 (N3555, N3253, N3488);
nand NAND2_1047 (N3556, N3256, N3490);
nand NAND2_1048 (N3557, N3259, N3492);
and AND2_1049 (N3558, N3453, N3091);
and AND2_1050 (N3559, N3450, N3088);
nand NAND2_1051 (N3563, N3262, N3501);
nand NAND2_1052 (N3564, N3265, N3503);
nand NAND2_1053 (N3565, N3268, N3505);
nand NAND2_1054 (N3566, N3271, N3507);
nand NAND2_1055 (N3567, N3274, N3509);
nand NAND2_1056 (N3568, N3277, N3511);
and AND2_1057 (N3569, N3459, N3113);
and AND2_1058 (N3570, N3456, N3110);
buf BUFF1_1059 (N3576, N3453);
buf BUFF1_1060 (N3579, N3450);
buf BUFF1_1061 (N3585, N3459);
buf BUFF1_1062 (N3588, N3456);
not NOT1_1063 (N3592, N3522);
nand NAND2_1064 (N3593, N3522, N3405);
not NOT1_1065 (N3594, N3525);
nand NAND2_1066 (N3595, N3525, N3406);
not NOT1_1067 (N3596, N3528);
nand NAND2_1068 (N3597, N3528, N2630);
nand NAND2_1069 (N3598, N3531, N2376);
not NOT1_1070 (N3599, N3531);
and AND2_1071 (N3600, N3551, N800);
nand NAND2_1072 (N3603, N3552, N3483);
nand NAND2_1073 (N3608, N3553, N3485);
nand NAND2_1074 (N3612, N3554, N3487);
nand NAND2_1075 (N3615, N3555, N3489);
nand NAND2_1076 (N3616, N3556, N3491);
nand NAND2_1077 (N3622, N3557, N3493);
not NOT1_1078 (N3629, N3534);
nand NAND2_1079 (N3630, N3534, N2645);
not NOT1_1080 (N3631, N3537);
nand NAND2_1081 (N3632, N3537, N2655);
nand NAND2_1082 (N3633, N3540, N2403);
not NOT1_1083 (N3634, N3540);
nand NAND2_1084 (N3635, N3563, N3502);
nand NAND2_1085 (N3640, N3564, N3504);
nand NAND2_1086 (N3644, N3565, N3506);
nand NAND2_1087 (N3647, N3566, N3508);
nand NAND2_1088 (N3648, N3567, N3510);
nand NAND2_1089 (N3654, N3568, N3512);
not NOT1_1090 (N3661, N3543);
nand NAND2_1091 (N3662, N3543, N2656);
nand NAND2_1092 (N3667, N3238, N3592);
nand NAND2_1093 (N3668, N3241, N3594);
nand NAND2_1094 (N3669, N2472, N3596);
nand NAND2_1095 (N3670, N2213, N3599);
buf BUFF1_1096 (dN3671, N3600);
not NOT1_1097 (N3691, N3576);
nand NAND2_1098 (N3692, N3576, N3494);
not NOT1_1099 (N3693, N3579);
nand NAND2_1100 (N3694, N3579, N3496);
nand NAND2_1101 (N3695, N2475, N3629);
nand NAND2_1102 (N3696, N2478, N3631);
nand NAND2_1103 (N3697, N2216, N3634);
not NOT1_1104 (N3716, N3585);
nand NAND2_1105 (N3717, N3585, N3513);
not NOT1_1106 (N3718, N3588);
nand NAND2_1107 (N3719, N3588, N3515);
nand NAND2_1108 (N3720, N2481, N3661);
nand NAND2_1109 (N3721, N3667, N3593);
nand NAND2_1110 (N3722, N3668, N3595);
nand NAND2_1111 (N3723, N3669, N3597);
nand NAND2_1112 (N3726, N3670, N3598);
not NOT1_1113 (N3727, N3600);
nand NAND2_1114 (N3728, N3364, N3691);
nand NAND2_1115 (N3729, N3367, N3693);
nand NAND2_1116 (N3730, N3695, N3630);
and AND4_1117 (N3731, N3608, N3615, N3612, N3603);
and AND2_1118 (N3732, N3603, N3293);
and AND3_1119 (N3733, N3608, N3603, N3295);
and AND4_1120 (N3734, N3612, N3603, N3296, N3608);
and AND2_1121 (N3735, N3616, N3301);
and AND3_1122 (N3736, N3622, N3616, N3558);
nand NAND2_1123 (N3737, N3696, N3632);
nand NAND2_1124 (N3740, N3697, N3633);
nand NAND2_1125 (N3741, N3394, N3716);
nand NAND2_1126 (N3742, N3397, N3718);
nand NAND2_1127 (N3743, N3720, N3662);
and AND4_1128 (N3744, N3640, N3647, N3644, N3635);
and AND2_1129 (N3745, N3635, N3306);
and AND3_1130 (N3746, N3640, N3635, N3308);
and AND4_1131 (N3747, N3644, N3635, N3309, N3640);
and AND2_1132 (N3748, N3648, N3314);
and AND3_1133 (N3749, N3654, N3648, N3569);
not NOT1_1134 (N3750, N3721);
and AND2_1135 (N3753, N3722, dN246);
nand NAND2_1136 (N3754, N3728, N3692);
nand NAND2_1137 (N3758, N3729, N3694);
not NOT1_1138 (N3761, N3731);
or OR4_1139 (N3762, N3291, N3732, N3733, N3734);
nand NAND2_1140 (N3767, N3741, N3717);
nand NAND2_1141 (N3771, N3742, N3719);
not NOT1_1142 (N3774, N3744);
or OR4_1143 (N3775, N3304, N3745, N3746, N3747);
and AND2_1144 (N3778, N3723, N3480);
and AND3_1145 (N3779, N3726, N3723, N3409);
or OR2_1146 (N3780, N2125, N3753);
and AND2_1147 (N3790, N3750, N800);
and AND2_1148 (N3793, N3737, N3500);
and AND3_1149 (N3794, N3740, N3737, N3428);
or OR3_1150 (N3802, N3479, N3778, N3779);
buf BUFF1_1151 (dN3803, N3780);
buf BUFF1_1152 (dN3804, N3780);
not NOT1_1153 (N3805, N3762);
and AND5_1154 (N3806, N3622, N3730, N3754, N3616, N3758);
and AND4_1155 (N3807, N3754, N3616, N3559, N3622);
and AND5_1156 (N3808, N3758, N3754, N3616, N3498, N3622);
buf BUFF1_1157 (dN3809, N3790);
or OR3_1158 (N3811, N3499, N3793, N3794);
not NOT1_1159 (N3812, N3775);
and AND5_1160 (N3813, N3654, N3743, N3767, N3648, N3771);
and AND4_1161 (N3814, N3767, N3648, N3570, N3654);
and AND5_1162 (N3815, N3771, N3767, N3648, N3517, N3654);
or OR5_1163 (N3816, N3299, N3735, N3736, N3807, N3808);
and AND2_1164 (N3817, N3806, N3802);
nand NAND2_1165 (N3818, N3805, N3761);
not NOT1_1166 (N3819, N3790);
or OR5_1167 (N3820, N3312, N3748, N3749, N3814, N3815);
and AND2_1168 (N3821, N3813, N3811);
nand NAND2_1169 (N3822, N3812, N3774);
or OR2_1170 (N3823, N3816, N3817);
and AND3_1171 (N3826, N3727, N3819, N2841);
or OR2_1172 (N3827, N3820, N3821);
not NOT1_1173 (N3834, N3823);
and AND2_1174 (N3835, N3818, N3823);
not NOT1_1175 (N3836, N3827);
and AND2_1176 (N3837, N3822, N3827);
and AND2_1177 (N3838, N3762, N3834);
and AND2_1178 (N3839, N3775, N3836);
or OR2_1179 (N3840, N3838, N3835);
or OR2_1180 (N3843, N3839, N3837);
buf BUFF1_1181 (dN3851, N3843);
nand NAND2_1182 (N3852, N3843, N3840);
and AND2_1183 (N3857, N3843, N3852);
and AND2_1184 (N3858, N3852, N3840);
or OR2_1185 (N3859, N3857, N3858);
not NOT1_1186 (N3864, N3859);
and AND2_1187 (N3869, N3859, N3864);
or OR2_1188 (N3870, N3869, N3864);
not NOT1_1189 (dN3875, N3870);
and AND3_1190 (N3876, N2826, N3028, N3870);
and AND3_1191 (N3877, N3826, N3876, N1591);
buf BUFF1_1192 (dN3881, N3877);
not NOT1_1193 (dN3882, N3877);
buf BUFF1_1194 (dN143_O, dN143_I);
buf BUFF1_1195 (dN144_O, dN144_I);
buf BUFF1_1196 (dN145_O, dN145_I);
buf BUFF1_1197 (dN146_O, dN146_I);
buf BUFF1_1198 (dN147_O, dN147_I);
buf BUFF1_1199 (dN148_O, dN148_I);
buf BUFF1_1200 (dN149_O, dN149_I);
buf BUFF1_1201 (dN150_O, dN150_I);
buf BUFF1_1202 (dN151_O, dN151_I);
buf BUFF1_1203 (dN152_O, dN152_I);
buf BUFF1_1204 (dN153_O, dN153_I);
buf BUFF1_1205 (dN154_O, dN154_I);
buf BUFF1_1206 (dN155_O, dN155_I);
buf BUFF1_1207 (dN156_O, dN156_I);
buf BUFF1_1208 (dN157_O, dN157_I);
buf BUFF1_1209 (dN158_O, dN158_I);
buf BUFF1_1210 (dN159_O, dN159_I);
buf BUFF1_1211 (dN160_O, dN160_I);
buf BUFF1_1212 (dN161_O, dN161_I);
buf BUFF1_1213 (dN162_O, dN162_I);
buf BUFF1_1214 (dN163_O, dN163_I);
buf BUFF1_1215 (dN164_O, dN164_I);
buf BUFF1_1216 (dN165_O, dN165_I);
buf BUFF1_1217 (dN166_O, dN166_I);
buf BUFF1_1218 (dN167_O, dN167_I);
buf BUFF1_1219 (dN168_O, dN168_I);
buf BUFF1_1220 (dN169_O, dN169_I);
buf BUFF1_1221 (dN170_O, dN170_I);
buf BUFF1_1222 (dN171_O, dN171_I);
buf BUFF1_1223 (dN172_O, dN172_I);
buf BUFF1_1224 (dN173_O, dN173_I);
buf BUFF1_1225 (dN174_O, dN174_I);
buf BUFF1_1226 (dN175_O, dN175_I);
buf BUFF1_1227 (dN176_O, dN176_I);
buf BUFF1_1228 (dN177_O, dN177_I);
buf BUFF1_1229 (dN178_O, dN178_I);
buf BUFF1_1230 (dN179_O, dN179_I);
buf BUFF1_1231 (dN180_O, dN180_I);
buf BUFF1_1232 (dN181_O, dN181_I);
buf BUFF1_1233 (dN182_O, dN182_I);
buf BUFF1_1234 (dN183_O, dN183_I);
buf BUFF1_1235 (dN184_O, dN184_I);
buf BUFF1_1236 (dN185_O, dN185_I);
buf BUFF1_1237 (dN186_O, dN186_I);
buf BUFF1_1238 (dN187_O, dN187_I);
buf BUFF1_1239 (dN188_O, dN188_I);
buf BUFF1_1240 (dN189_O, dN189_I);
buf BUFF1_1241 (dN190_O, dN190_I);
buf BUFF1_1242 (dN191_O, dN191_I);
buf BUFF1_1243 (dN192_O, dN192_I);
buf BUFF1_1244 (dN193_O, dN193_I);
buf BUFF1_1245 (dN194_O, dN194_I);
buf BUFF1_1246 (dN195_O, dN195_I);
buf BUFF1_1247 (dN196_O, dN196_I);
buf BUFF1_1248 (dN197_O, dN197_I);
buf BUFF1_1249 (dN198_O, dN198_I);
buf BUFF1_1250 (dN199_O, dN199_I);
buf BUFF1_1251 (dN200_O, dN200_I);
buf BUFF1_1252 (dN201_O, dN201_I);
buf BUFF1_1253 (dN202_O, dN202_I);
buf BUFF1_1254 (dN203_O, dN203_I);
buf BUFF1_1255 (dN204_O, dN204_I);
buf BUFF1_1256 (dN205_O, dN205_I);
buf BUFF1_1257 (dN206_O, dN206_I);
buf BUFF1_1258 (dN207_O, dN207_I);
buf BUFF1_1259 (dN208_O, dN208_I);
buf BUFF1_1260 (dN209_O, dN209_I);
buf BUFF1_1261 (dN210_O, dN210_I);
buf BUFF1_1262 (dN211_O, dN211_I);
buf BUFF1_1263 (dN212_O, dN212_I);
buf BUFF1_1264 (dN213_O, dN213_I);
buf BUFF1_1265 (dN214_O, dN214_I);
buf BUFF1_1266 (dN215_O, dN215_I);
buf BUFF1_1267 (dN216_O, dN216_I);
buf BUFF1_1268 (dN217_O, dN217_I);
buf BUFF1_1269 (dN218_O, dN218_I);

// D Flip-Flops in front of input	
dff a1 (dN1, N1, clk);
dff a2 (dN2, N2, clk);
dff a3 (dN3, N3, clk);
dff a4 (dN4, N4, clk);
dff a5 (dN5, N5, clk);
dff a6 (dN6, N6, clk);
dff a7 (dN7, N7, clk);
dff a8 (dN8, N8, clk);
dff a9 (dN11, N11, clk);
dff a10 (dN14, N14, clk);
dff a11 (dN15, N15, clk);
dff a12 (dN16, N16, clk);
dff a13 (dN19, N19, clk);
dff a14 (dN20, N20, clk);
dff a15 (dN21, N21, clk);
dff a16 (dN22, N22, clk);
dff a17 (dN23, N23, clk);
dff a18 (dN24, N24, clk);
dff a19 (dN25, N25, clk);
dff a20 (dN26, N26, clk);
dff a21 (dN27, N27, clk);
dff a22 (dN28, N28, clk);
dff a23 (dN29, N29, clk);
dff a24 (dN32, N32, clk);
dff a25 (dN33, N33, clk);
dff a26 (dN34, N34, clk);
dff a27 (dN35, N35, clk);
dff a28 (dN36, N36, clk);
dff a29 (dN37, N37, clk);
dff a30 (dN40, N40, clk);
dff a31 (dN43, N43, clk);
dff a32 (dN44, N44, clk);
dff a33 (dN47, N47, clk);
dff a34 (dN48, N48, clk);
dff a35 (dN49, N49, clk);
dff a36 (dN50, N50, clk);
dff a37 (dN51, N51, clk);
dff a38 (dN52, N52, clk);
dff a39 (dN53, N53, clk);
dff a40 (dN54, N54, clk);
dff a41 (dN55, N55, clk);
dff a42 (dN56, N56, clk);
dff a43 (dN57, N57, clk);
dff a44 (dN60, N60, clk);
dff a45 (dN61, N61, clk);
dff a46 (dN62, N62, clk);
dff a47 (dN63, N63, clk);
dff a48 (dN64, N64, clk);
dff a49 (dN65, N65, clk);
dff a50 (dN66, N66, clk);
dff a51 (dN67, N67, clk);
dff a52 (dN68, N68, clk);
dff a53 (dN69, N69, clk);
dff a54 (dN72, N72, clk);
dff a55 (dN73, N73, clk);
dff a56 (dN74, N74, clk);
dff a57 (dN75, N75, clk);
dff a58 (dN76, N76, clk);
dff a59 (dN77, N77, clk);
dff a60 (dN78, N78, clk);
dff a61 (dN79, N79, clk);
dff a62 (dN80, N80, clk);
dff a63 (dN81, N81, clk);
dff a64 (dN82, N82, clk);
dff a65 (dN85, N85, clk);
dff a66 (dN86, N86, clk);
dff a67 (dN87, N87, clk);
dff a68 (dN88, N88, clk);
dff a69 (dN89, N89, clk);
dff a70 (dN90, N90, clk);
dff a71 (dN91, N91, clk);
dff a72 (dN92, N92, clk);
dff a73 (dN93, N93, clk);
dff a74 (dN94, N94, clk);
dff a75 (dN95, N95, clk);
dff a76 (dN96, N96, clk);
dff a77 (dN99, N99, clk);
dff a78 (dN100, N100, clk);
dff a79 (dN101, N101, clk);
dff a80 (dN102, N102, clk);
dff a81 (dN103, N103, clk);
dff a82 (dN104, N104, clk);
dff a83 (dN105, N105, clk);
dff a84 (dN106, N106, clk);
dff a85 (dN107, N107, clk);
dff a86 (dN108, N108, clk);
dff a87 (dN111, N111, clk);
dff a88 (dN112, N112, clk);
dff a89 (dN113, N113, clk);
dff a90 (dN114, N114, clk);
dff a91 (dN115, N115, clk);
dff a92 (dN116, N116, clk);
dff a93 (dN117, N117, clk);
dff a94 (dN118, N118, clk);
dff a95 (dN119, N119, clk);
dff a96 (dN120, N120, clk);
dff a97 (dN123, N123, clk);
dff a98 (dN124, N124, clk);
dff a99 (dN125, N125, clk);
dff a100 (dN126, N126, clk);
dff a101 (dN127, N127, clk);
dff a102 (dN128, N128, clk);
dff a103 (dN129, N129, clk);
dff a104 (dN130, N130, clk);
dff a105 (dN131, N131, clk);
dff a106 (dN132, N132, clk);
dff a107 (dN135, N135, clk);
dff a108 (dN136, N136, clk);
dff a109 (dN137, N137, clk);
dff a110 (dN138, N138, clk);
dff a111 (dN139, N139, clk);
dff a112 (dN140, N140, clk);
dff a113 (dN141, N141, clk);
dff a114 (dN142, N142, clk);
dff a115 (dN219, N219, clk);
dff a116 (dN224, N224, clk);
dff a117 (dN227, N227, clk);
dff a118 (dN230, N230, clk);
dff a119 (dN231, N231, clk);
dff a120 (dN234, N234, clk);
dff a121 (dN237, N237, clk);
dff a122 (dN241, N241, clk);
dff a123 (dN246, N246, clk);
dff a124 (dN253, N253, clk);
dff a125 (dN256, N256, clk);
dff a126 (dN259, N259, clk);
dff a127 (dN262, N262, clk);
dff a128 (dN263, N263, clk);
dff a129 (dN266, N266, clk);
dff a130 (dN269, N269, clk);
dff a131 (dN272, N272, clk);
dff a132 (dN275, N275, clk);
dff a133 (dN278, N278, clk);
dff a134 (dN281, N281, clk);
dff a135 (dN284, N284, clk);
dff a136 (dN287, N287, clk);
dff a137 (dN290, N290, clk);
dff a138 (dN294, N294, clk);
dff a139 (dN297, N297, clk);
dff a140 (dN301, N301, clk);
dff a141 (dN305, N305, clk);
dff a142 (dN309, N309, clk);
dff a143 (dN313, N313, clk);
dff a144 (dN316, N316, clk);
dff a145 (dN319, N319, clk);
dff a146 (dN322, N322, clk);
dff a147 (dN325, N325, clk);
dff a148 (dN328, N328, clk);
dff a149 (dN331, N331, clk);
dff a150 (dN334, N334, clk);
dff a151 (dN337, N337, clk);
dff a152 (dN340, N340, clk);
dff a153 (dN343, N343, clk);
dff a154 (dN346, N346, clk);
dff a155 (dN349, N349, clk);
dff a156 (dN352, N352, clk);
dff a157 (dN355, N355, clk);
dff a158 (dN143_I, N143_I, clk);
dff a159 (dN144_I, N144_I, clk);
dff a160 (dN145_I, N145_I, clk);
dff a161 (dN146_I, N146_I, clk);
dff a162 (dN147_I, N147_I, clk);
dff a163 (dN148_I, N148_I, clk);
dff a164 (dN149_I, N149_I, clk);
dff a165 (dN150_I, N150_I, clk);
dff a166 (dN151_I, N151_I, clk);
dff a167 (dN152_I, N152_I, clk);
dff a168 (dN153_I, N153_I, clk);
dff a169 (dN154_I, N154_I, clk);
dff a170 (dN155_I, N155_I, clk);
dff a171 (dN156_I, N156_I, clk);
dff a172 (dN157_I, N157_I, clk);
dff a173 (dN158_I, N158_I, clk);
dff a174 (dN159_I, N159_I, clk);
dff a175 (dN160_I, N160_I, clk);
dff a176 (dN161_I, N161_I, clk);
dff a177 (dN162_I, N162_I, clk);
dff a178 (dN163_I, N163_I, clk);
dff a179 (dN164_I, N164_I, clk);
dff a180 (dN165_I, N165_I, clk);
dff a181 (dN166_I, N166_I, clk);
dff a182 (dN167_I, N167_I, clk);
dff a183 (dN168_I, N168_I, clk);
dff a184 (dN169_I, N169_I, clk);
dff a185 (dN170_I, N170_I, clk);
dff a186 (dN171_I, N171_I, clk);
dff a187 (dN172_I, N172_I, clk);
dff a188 (dN173_I, N173_I, clk);
dff a189 (dN174_I, N174_I, clk);
dff a190 (dN175_I, N175_I, clk);
dff a191 (dN176_I, N176_I, clk);
dff a192 (dN177_I, N177_I, clk);
dff a193 (dN178_I, N178_I, clk);
dff a194 (dN179_I, N179_I, clk);
dff a195 (dN180_I, N180_I, clk);
dff a196 (dN181_I, N181_I, clk);
dff a197 (dN182_I, N182_I, clk);
dff a198 (dN183_I, N183_I, clk);
dff a199 (dN184_I, N184_I, clk);
dff a200 (dN185_I, N185_I, clk);
dff a201 (dN186_I, N186_I, clk);
dff a202 (dN187_I, N187_I, clk);
dff a203 (dN188_I, N188_I, clk);
dff a204 (dN189_I, N189_I, clk);
dff a205 (dN190_I, N190_I, clk);
dff a206 (dN191_I, N191_I, clk);
dff a207 (dN192_I, N192_I, clk);
dff a208 (dN193_I, N193_I, clk);
dff a209 (dN194_I, N194_I, clk);
dff a210 (dN195_I, N195_I, clk);
dff a211 (dN196_I, N196_I, clk);
dff a212 (dN197_I, N197_I, clk);
dff a213 (dN198_I, N198_I, clk);
dff a214 (dN199_I, N199_I, clk);
dff a215 (dN200_I, N200_I, clk);
dff a216 (dN201_I, N201_I, clk);
dff a217 (dN202_I, N202_I, clk);
dff a218 (dN203_I, N203_I, clk);
dff a219 (dN204_I, N204_I, clk);
dff a220 (dN205_I, N205_I, clk);
dff a221 (dN206_I, N206_I, clk);
dff a222 (dN207_I, N207_I, clk);
dff a223 (dN208_I, N208_I, clk);
dff a224 (dN209_I, N209_I, clk);
dff a225 (dN210_I, N210_I, clk);
dff a226 (dN211_I, N211_I, clk);
dff a227 (dN212_I, N212_I, clk);
dff a228 (dN213_I, N213_I, clk);
dff a229 (dN214_I, N214_I, clk);
dff a230 (dN215_I, N215_I, clk);
dff a231 (dN216_I, N216_I, clk);
dff a232 (dN217_I, N217_I, clk);
dff a233 (dN218_I, N218_I, clk);
	
	
// D Flip-Flops after output
dff b1 (N398, dN398, clk);
dff b2 (N400, dN400, clk);
dff b3 (N401, dN401, clk);
dff b4 (N419, dN419, clk);
dff b5 (N420, dN420, clk);
dff b6 (N456, dN456, clk);
dff b7 (N457, dN457, clk);
dff b8 (N458, dN458, clk);
dff b9 (N487, dN487, clk);
dff b10 (N488, dN488, clk);
dff b11 (N489, dN489, clk);
dff b12 (N490, dN490, clk);
dff b13 (N491, dN491, clk);
dff b14 (N492, dN492, clk);
dff b15 (N493, dN493, clk);
dff b16 (N494, dN494, clk);
dff b17 (N792, dN792, clk);
dff b18 (N799, dN799, clk);
dff b19 (N805, dN805, clk);
dff b20 (N1026, dN1026, clk);
dff b21 (N1028, dN1028, clk);
dff b22 (N1029, dN1029, clk);
dff b23 (N1269, dN1269, clk);
dff b24 (N1277, dN1277, clk);
dff b25 (N1448, dN1448, clk);
dff b26 (N1726, dN1726, clk);
dff b27 (N1816, dN1816, clk);
dff b28 (N1817, dN1817, clk);
dff b29 (N1818, dN1818, clk);
dff b30 (N1819, dN1819, clk);
dff b31 (N1820, dN1820, clk);
dff b32 (N1821, dN1821, clk);
dff b33 (N1969, dN1969, clk);
dff b34 (N1970, dN1970, clk);
dff b35 (N1971, dN1971, clk);
dff b36 (N2010, dN2010, clk);
dff b37 (N2012, dN2012, clk);
dff b38 (N2014, dN2014, clk);
dff b39 (N2016, dN2016, clk);
dff b40 (N2018, dN2018, clk);
dff b41 (N2020, dN2020, clk);
dff b42 (N2022, dN2022, clk);
dff b43 (N2387, dN2387, clk);
dff b44 (N2388, dN2388, clk);
dff b45 (N2389, dN2389, clk);
dff b46 (N2390, dN2390, clk);
dff b47 (N2496, dN2496, clk);
dff b48 (N2643, dN2643, clk);
dff b49 (N2644, dN2644, clk);
dff b50 (N2891, dN2891, clk);
dff b51 (N2925, dN2925, clk);
dff b52 (N2970, dN2970, clk);
dff b53 (N2971, dN2971, clk);
dff b54 (N3038, dN3038, clk);
dff b55 (N3079, dN3079, clk);
dff b56 (N3546, dN3546, clk);
dff b57 (N3671, dN3671, clk);
dff b58 (N3803, dN3803, clk);
dff b59 (N3804, dN3804, clk);
dff b60 (N3809, dN3809, clk);
dff b61 (N3851, dN3851, clk);
dff b62 (N3875, dN3875, clk);
dff b63 (N3881, dN3881, clk);
dff b64 (N3882, dN3882, clk);
dff b65 (N143_O, dN143_O, clk);
dff b66 (N144_O, dN144_O, clk);
dff b67 (N145_O, dN145_O, clk);
dff b68 (N146_O, dN146_O, clk);
dff b69 (N147_O, dN147_O, clk);
dff b70 (N148_O, dN148_O, clk);
dff b71 (N149_O, dN149_O, clk);
dff b72 (N150_O, dN150_O, clk);
dff b73 (N151_O, dN151_O, clk);
dff b74 (N152_O, dN152_O, clk);
dff b75 (N153_O, dN153_O, clk);
dff b76 (N154_O, dN154_O, clk);
dff b77 (N155_O, dN155_O, clk);
dff b78 (N156_O, dN156_O, clk);
dff b79 (N157_O, dN157_O, clk);
dff b80 (N158_O, dN158_O, clk);
dff b81 (N159_O, dN159_O, clk);
dff b82 (N160_O, dN160_O, clk);
dff b83 (N161_O, dN161_O, clk);
dff b84 (N162_O, dN162_O, clk);
dff b85 (N163_O, dN163_O, clk);
dff b86 (N164_O, dN164_O, clk);
dff b87 (N165_O, dN165_O, clk);
dff b88 (N166_O, dN166_O, clk);
dff b89 (N167_O, dN167_O, clk);
dff b90 (N168_O, dN168_O, clk);
dff b91 (N169_O, dN169_O, clk);
dff b92 (N170_O, dN170_O, clk);
dff b93 (N171_O, dN171_O, clk);
dff b94 (N172_O, dN172_O, clk);
dff b95 (N173_O, dN173_O, clk);
dff b96 (N174_O, dN174_O, clk);
dff b97 (N175_O, dN175_O, clk);
dff b98 (N176_O, dN176_O, clk);
dff b99 (N177_O, dN177_O, clk);
dff b100 (N178_O, dN178_O, clk);
dff b101 (N179_O, dN179_O, clk);
dff b102 (N180_O, dN180_O, clk);
dff b103 (N181_O, dN181_O, clk);
dff b104 (N182_O, dN182_O, clk);
dff b105 (N183_O, dN183_O, clk);
dff b106 (N184_O, dN184_O, clk);
dff b107 (N185_O, dN185_O, clk);
dff b108 (N186_O, dN186_O, clk);
dff b109 (N187_O, dN187_O, clk);
dff b110 (N188_O, dN188_O, clk);
dff b111 (N189_O, dN189_O, clk);
dff b112 (N190_O, dN190_O, clk);
dff b113 (N191_O, dN191_O, clk);
dff b114 (N192_O, dN192_O, clk);
dff b115 (N193_O, dN193_O, clk);
dff b116 (N194_O, dN194_O, clk);
dff b117 (N195_O, dN195_O, clk);
dff b118 (N196_O, dN196_O, clk);
dff b119 (N197_O, dN197_O, clk);
dff b120 (N198_O, dN198_O, clk);
dff b121 (N199_O, dN199_O, clk);
dff b122 (N200_O, dN200_O, clk);
dff b123 (N201_O, dN201_O, clk);
dff b124 (N202_O, dN202_O, clk);
dff b125 (N203_O, dN203_O, clk);
dff b126 (N204_O, dN204_O, clk);
dff b127 (N205_O, dN205_O, clk);
dff b128 (N206_O, dN206_O, clk);
dff b129 (N207_O, dN207_O, clk);
dff b130 (N208_O, dN208_O, clk);
dff b131 (N209_O, dN209_O, clk);
dff b132 (N210_O, dN210_O, clk);
dff b133 (N211_O, dN211_O, clk);
dff b134 (N212_O, dN212_O, clk);
dff b135 (N213_O, dN213_O, clk);
dff b136 (N214_O, dN214_O, clk);
dff b137 (N215_O, dN215_O, clk);
dff b138 (N216_O, dN216_O, clk);
dff b139 (N217_O, dN217_O, clk);
dff b140 (N218_O, dN218_O, clk);

endmodule

module dff(q, d, clk);
	input  d, clk;
	output reg q;

always @ (posedge clk)
	q <= d;
	
endmodule

//------------------------------------------------------------------------------------------------------------------------------------------------------
//---------------------------------------------------------------------------------------------------------------------------------------------------
`timescale 1ns/ 1ps

module Testbench_benchmarkc2670();

reg clk, en, N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22, N23, N24, N25, N26,  N27, N28, N29, N32, N33, N34, N35, N36, N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54,  N55, N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76, N77, N78,  N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N99, N100, N101, N102,  N103, N104, N105, N106, N107, N108, N111, N112, N113, N114,  N115, N116, N117, N118, N119, N120, N123, N124, N125, N126,  N127, N128, N129, N130, N131, N132, N135, N136, N137, N138,  N139, N140, N141, N142, N219, N224, N227, N230, N231, N234,  N237, N241, N246, N253, N256, N259, N262, N263, N266, N269,  N272, N275, N278, N281, N284, N287, N290, N294, N297, N301,  N305, N309, N313, N316, N319, N322, N325, N328, N331, N334,  N337, N340, N343, N346, N349, N352, N355, N143_I, N144_I, N145_I,  N146_I, N147_I, N148_I, N149_I, N150_I, N151_I, N152_I, N153_I, N154_I, N155_I,  N156_I, N157_I, N158_I, N159_I, N160_I, N161_I, N162_I, N163_I, N164_I, N165_I,  N166_I, N167_I, N168_I, N169_I, N170_I, N171_I, N172_I, N173_I, N174_I, N175_I,  N176_I, N177_I, N178_I, N179_I, N180_I, N181_I, N182_I, N183_I, N184_I, N185_I,  N186_I, N187_I, N188_I, N189_I, N190_I, N191_I, N192_I, N193_I, N194_I, N195_I,  N196_I, N197_I, N198_I, N199_I, N200_I, N201_I, N202_I, N203_I, N204_I, N205_I,  N206_I, N207_I, N208_I, N209_I, N210_I, N211_I, N212_I, N213_I, N214_I, N215_I,  N216_I, N217_I, N218_I;

wire N398, N400, N401, N419, N420, N456, N457, N458, N487, N488, N489, N490, N491, N492, N493, N494, N792, N799, N805, N1026, N1028, N1029, N1269, N1277, N1448, N1726, N1816, N1817, N1818, N1819, N1820, N1821, N1969, N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022, N2387, N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925, N2970, N2971, N3038, N3079, N3546, N3671, N3803, N3804, N3809, N3851, N3875, N3881, N3882, N143_O, N144_O, N145_O, N146_O, N147_O, N148_O, N149_O, N150_O, N151_O, N152_O, N153_O, N154_O, N155_O, N156_O, N157_O, N158_O, N159_O, N160_O, N161_O, N162_O, N163_O, N164_O, N165_O, N166_O, N167_O, N168_O, N169_O, N170_O, N171_O, N172_O, N173_O, N174_O, N175_O, N176_O, N177_O, N178_O, N179_O, N180_O, N181_O, N182_O, N183_O, N184_O, N185_O, N186_O, N187_O, N188_O, N189_O, N190_O, N191_O, N192_O, N193_O, N194_O, N195_O, N196_O, N197_O, N198_O, N199_O, N200_O, N201_O, N202_O, N203_O, N204_O, N205_O, N206_O, N207_O, N208_O, N209_O, N210_O, N211_O, N212_O, N213_O, N214_O, N215_O, N216_O, N217_O, N218_O;

 //instantiation
c2670 dut(
//input port mapping
	.clk(clk),
	.en(en),
	.N1(N1),
	.N2(N2),
	.N3(N3),
	.N4(N4),
	.N5(N5),
	.N6(N6),
	.N7(N7),
	.N8(N8),
	.N11(N11),
	.N14(N14),
	.N15(N15),
	.N16(N16),
	.N19(N19),
	.N20(N20),
	.N21(N21),
	.N22(N22),
	.N23(N23),
	.N24(N24),
	.N25(N25),
	.N26(N26),
	.N27(N27),
	.N28(N28),
	.N29(N29),
	.N32(N32),
	.N33(N33),
	.N34(N34),
	.N35(N35),
	.N36(N36),
	.N37(N37),
	.N40(N40),
	.N43(N43),
	.N44(N44),
	.N47(N47),
	.N48(N48),
	.N49(N49),
	.N50(N50),
	.N51(N51),
	.N52(N52),
	.N53(N53),
	.N54(N54),
	.N55(N55),
	.N56(N56),
	.N57(N57),
	.N60(N60),
	.N61(N61),
	.N62(N62),
	.N63(N63),
	.N64(N64),
	.N65(N65),
	.N66(N66),
	.N67(N67),
	.N68(N68),
	.N69(N69),
	.N72(N72),
	.N73(N73),
	.N74(N74),
	.N75(N75),
	.N76(N76),
	.N77(N77),
	.N78(N78),
	.N79(N79),
	.N80(N80),
	.N81(N81),
	.N82(N82),
	.N85(N85),
	.N86(N86),
	.N87(N87),
	.N88(N88),
	.N89(N89),
	.N90(N90),
	.N91(N91),
	.N92(N92),
	.N93(N93),
	.N94(N94),
	.N95(N95),
	.N96(N96),
	.N99(N99),
	.N100(N100),
	.N101(N101),
	.N102(N102),
	.N103(N103),
	.N104(N104),
	.N105(N105),
	.N106(N106),
	.N107(N107),
	.N108(N108),
	.N111(N111),
	.N112(N112),
	.N113(N113),
	.N114(N114),
	.N115(N115),
	.N116(N116),
	.N117(N117),
	.N118(N118),
	.N119(N119),
	.N120(N120),
	.N123(N123),
	.N124(N124),
	.N125(N125),
	.N126(N126),
	.N127(N127),
	.N128(N128),
	.N129(N129),
	.N130(N130),
	.N131(N131),
	.N132(N132),
	.N135(N135),
	.N136(N136),
	.N137(N137),
	.N138(N138),
	.N139(N139),
	.N140(N140),
	.N141(N141),
	.N142(N142),
	.N219(N219),
	.N224(N224),
	.N227(N227),
	.N230(N230),
	.N231(N231),
	.N234(N234),
	.N237(N237),
	.N241(N241),
	.N246(N246),
	.N253(N253),
	.N256(N256),
	.N259(N259),
	.N262(N262),
	.N263(N263),
	.N266(N266),
	.N269(N269),
	.N272(N272),
	.N275(N275),
	.N278(N278),
	.N281(N281),
	.N284(N284),
	.N287(N287),
	.N290(N290),
	.N294(N294),
	.N297(N297),
	.N301(N301),
	.N305(N305),
	.N309(N309),
	.N313(N313),
	.N316(N316),
	.N319(N319),
	.N322(N322),
	.N325(N325),
	.N328(N328),
	.N331(N331),
	.N334(N334),
	.N337(N337),
	.N340(N340),
	.N343(N343),
	.N346(N346),
	.N349(N349),
	.N352(N352),
	.N355(N355),
	.N143_I(N143_I),
	.N144_I(N144_I),
	.N145_I(N145_I),
	.N146_I(N146_I),
	.N147_I(N147_I),
	.N148_I(N148_I),
	.N149_I(N149_I),
	.N150_I(N150_I),
	.N151_I(N151_I),
	.N152_I(N152_I),
	.N153_I(N153_I),
	.N154_I(N154_I),
	.N155_I(N155_I),
	.N156_I(N156_I),
	.N157_I(N157_I),
	.N158_I(N158_I),
	.N159_I(N159_I),
	.N160_I(N160_I),
	.N161_I(N161_I),
	.N162_I(N162_I),
	.N163_I(N163_I),
	.N164_I(N164_I),
	.N165_I(N165_I),
	.N166_I(N166_I),
	.N167_I(N167_I),
	.N168_I(N168_I),
	.N169_I(N169_I),
	.N170_I(N170_I),
	.N171_I(N171_I),
	.N172_I(N172_I),
	.N173_I(N173_I),
	.N174_I(N174_I),
	.N175_I(N175_I),
	.N176_I(N176_I),
	.N177_I(N177_I),
	.N178_I(N178_I),
	.N179_I(N179_I),
	.N180_I(N180_I),
	.N181_I(N181_I),
	.N182_I(N182_I),
	.N183_I(N183_I),
	.N184_I(N184_I),
	.N185_I(N185_I),
	.N186_I(N186_I),
	.N187_I(N187_I),
	.N188_I(N188_I),
	.N189_I(N189_I),
	.N190_I(N190_I),
	.N191_I(N191_I),
	.N192_I(N192_I),
	.N193_I(N193_I),
	.N194_I(N194_I),
	.N195_I(N195_I),
	.N196_I(N196_I),
	.N197_I(N197_I),
	.N198_I(N198_I),
	.N199_I(N199_I),
	.N200_I(N200_I),
	.N201_I(N201_I),
	.N202_I(N202_I),
	.N203_I(N203_I),
	.N204_I(N204_I),
	.N205_I(N205_I),
	.N206_I(N206_I),
	.N207_I(N207_I),
	.N208_I(N208_I),
	.N209_I(N209_I),
	.N210_I(N210_I),
	.N211_I(N211_I),
	.N212_I(N212_I),
	.N213_I(N213_I),
	.N214_I(N214_I),
	.N215_I(N215_I),
	.N216_I(N216_I),
	.N217_I(N217_I),
	.N218_I(N218_I),
	
//output port mapping	
	.N398(N398),
	.N400(N400),
	.N401(N401),
	.N419(N419),
	.N420(N420),
	.N456(N456),
	.N457(N457),
	.N458(N458),
	.N487(N487),
	.N488(N488),
	.N489(N489),
	.N490(N490),
	.N491(N491),
	.N492(N492),
	.N493(N493),
	.N494(N494),
	.N792(N792),
	.N799(N799),
	.N805(N805),
	.N1026(N1026),
	.N1028(N1028),
	.N1029(N1029),
	.N1269(N1269),
	.N1277(N1277),
	.N1448(N1448),
	.N1726(N1726),
	.N1816(N1816),
	.N1817(N1817),
	.N1818(N1818),
	.N1819(N1819),
	.N1820(N1820),
	.N1821(N1821),
	.N1969(N1969),
	.N1970(N1970),
	.N1971(N1971),
	.N2010(N2010),
	.N2012(N2012),
	.N2014(N2014),
	.N2016(N2016),
	.N2018(N2018),
	.N2020(N2020),
	.N2022(N2022),
	.N2387(N2387),
	.N2388(N2388),
	.N2389(N2389),
	.N2390(N2390),
	.N2496(N2496),
	.N2643(N2643),
	.N2644(N2644),
	.N2891(N2891),
	.N2925(N2925),
	.N2970(N2970),
	.N2971(N2971),
	.N3038(N3038),
	.N3079(N3079),
	.N3546(N3546),
	.N3671(N3671),
	.N3803(N3803),
	.N3804(N3804),
	.N3809(N3809),
	.N3851(N3851),
	.N3875(N3875),
	.N3881(N3881),
	.N3882(N3882),
	.N143_O(N143_O),
	.N144_O(N144_O),
	.N145_O(N145_O),
	.N146_O(N146_O),
	.N147_O(N147_O),
	.N148_O(N148_O),
	.N149_O(N149_O),
	.N150_O(N150_O),
	.N151_O(N151_O),
	.N152_O(N152_O),
	.N153_O(N153_O),
	.N154_O(N154_O),
	.N155_O(N155_O),
	.N156_O(N156_O),
	.N157_O(N157_O),
	.N158_O(N158_O),
	.N159_O(N159_O),
	.N160_O(N160_O),
	.N161_O(N161_O),
	.N162_O(N162_O),
	.N163_O(N163_O),
	.N164_O(N164_O),
	.N165_O(N165_O),
	.N166_O(N166_O),
	.N167_O(N167_O),
	.N168_O(N168_O),
	.N169_O(N169_O),
	.N170_O(N170_O),
	.N171_O(N171_O),
	.N172_O(N172_O),
	.N173_O(N173_O),
	.N174_O(N174_O),
	.N175_O(N175_O),
	.N176_O(N176_O),
	.N177_O(N177_O),
	.N178_O(N178_O),
	.N179_O(N179_O),
	.N180_O(N180_O),
	.N181_O(N181_O),
	.N182_O(N182_O),
	.N183_O(N183_O),
	.N184_O(N184_O),
	.N185_O(N185_O),
	.N186_O(N186_O),
	.N187_O(N187_O),
	.N188_O(N188_O),
	.N189_O(N189_O),
	.N190_O(N190_O),
	.N191_O(N191_O),
	.N192_O(N192_O),
	.N193_O(N193_O),
	.N194_O(N194_O),
	.N195_O(N195_O),
	.N196_O(N196_O),
	.N197_O(N197_O),
	.N198_O(N198_O),
	.N199_O(N199_O),
	.N200_O(N200_O),
	.N201_O(N201_O),
	.N202_O(N202_O),
	.N203_O(N203_O),
	.N204_O(N204_O),
	.N205_O(N205_O),
	.N206_O(N206_O),
	.N207_O(N207_O),
	.N208_O(N208_O),
	.N209_O(N209_O),
	.N210_O(N210_O),
	.N211_O(N211_O),
	.N212_O(N212_O),
	.N213_O(N213_O),
	.N214_O(N214_O),
	.N215_O(N215_O),
	.N216_O(N216_O),
	.N217_O(N217_O),
	.N218_O(N218_O)
);
   

initial begin
	clk=0; en = 0; 
    N1=clk; N2=clk; N3=clk; N4=clk; N5=clk; N6=clk; N7=clk; N8=clk; N11=clk; N14=clk; N15=clk; N16=clk; N19=clk; N20=clk; N21=clk; N22=clk; N23=clk; N24=clk; N25=clk; N26=clk; N27=clk; N28=clk; 
	N29=clk; N32=clk; N33=clk; N34=clk; N35=clk; N36=clk; N37=clk; N40=clk; N43=clk; N44=clk; N47=clk; N48=clk; N49=clk; N50=clk; N51=clk; N52=clk; N53=clk; N54=clk; N55=clk; N56=clk; N57=clk; 
	N60=clk; N61=clk; N62=clk; N63=clk; N64=clk; N65=clk; N66=clk; N67=clk; N68=clk; N69=clk; N72=clk; N73=clk; N74=clk; N75=clk; N76=clk; N77=clk; N78=clk;  N79=clk; N80=clk; N81=clk; N82=clk; 
	N85=clk; N86=clk; N87=clk; N88=clk; N89=clk; N90=clk; N91=clk; N92=clk; N93=clk; N94=clk; N95=clk; N96=clk; N99=clk; N100=clk; N101=clk; N102=clk; N103=clk; N104=clk; N105=clk; N106=clk; 
	N107=clk; N108=clk; N111=clk; N112=clk; N113=clk; N114=clk; N115=clk; N116=clk; N117=clk; N118=clk; N119=clk; N120=clk; N123=clk; N124=clk; N125=clk; N126=clk; N127=clk; N128=clk; 
	N129=clk; N130=clk; N131=clk; N132=clk; N135=clk; N136=clk; N137=clk; N138=clk; N139=clk; N140=clk; N141=clk; N142=clk; N219=clk; N224=clk; N227=clk; N230=clk; N231=clk; N234=clk;  
	N237=clk; N241=clk; N246=clk; N253=clk; N256=clk; N259=clk; N262=clk; N263=clk; N266=clk; N269=clk; N272=clk; N275=clk; N278=clk; N281=clk; N284=clk; N287=clk; N290=clk; N294=clk; 
	N297=clk; N301=clk; N305=clk; N309=clk; N313=clk; N316=clk; N319=clk; N322=clk; N325=clk; N328=clk; N331=clk; N334=clk;  N337=clk; N340=clk; N343=clk; N346=clk; N349=clk; N352=clk; 
	N355=clk; N143_I=clk; N144_I=clk; N145_I=clk; N146_I=clk; N147_I=clk; N148_I=clk; N149_I=clk; N150_I=clk; N151_I=clk; N152_I=clk; N153_I=clk; N154_I=clk; N155_I=clk;  
	N156_I=clk; N157_I=clk; N158_I=clk; N159_I=clk; N160_I=clk; N161_I=clk; N162_I=clk; N163_I=clk; N164_I=clk; N165_I=clk; N166_I=clk; N167_I=clk; N168_I=clk; N169_I=clk; 
	N170_I=clk; N171_I=clk; N172_I=clk; N173_I=clk; N174_I=clk; N175_I=clk; N176_I=clk; N177_I=clk; N178_I=clk; N179_I=clk; N180_I=clk; N181_I=clk; N182_I=clk; N183_I=clk; 
	N184_I=clk; N185_I=clk; N186_I=clk; N187_I=clk; N188_I=clk; N189_I=clk; N190_I=clk; N191_I=clk; N192_I=clk; N193_I=clk; N194_I=clk; N195_I=clk; N196_I=clk; N197_I=clk; 
	N198_I=clk; N199_I=clk; N200_I=clk; N201_I=clk; N202_I=clk; N203_I=clk; N204_I=clk;  
	N205_I=clk;  N206_I=clk; N207_I=clk; N208_I=clk; N209_I=clk; N210_I=clk; N211_I=clk; N212_I=clk; N213_I=clk; N214_I=clk; N215_I=clk;  N216_I=clk; N217_I=clk; N218_I=clk;
	//$dumpfile ("c2670.vcd"); 
	//$dumpvars(0,Testbench_benchmarkc2670);

end

	always @ (posedge clk)
		$display("%3d,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b,%1b",$time,N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,N216_I,N217_I,N218_I,en,N398,N400,N401,N419,N420,N456,N457,N458,N487,N488,N489,N490,N491,N492,N493,N494,N792,N799,N805,N1026,N1028,N1029,N1269,N1277,N1448,N1726,N1816,N1817,N1818,N1819,N1820,N1821,N1969,N1970,N1971,N2010,N2012,N2014,N2016,N2018,N2020,N2022,N2387,N2388,N2389,N2390,N2496,N2643,N2644,N2891,N2925,N2970,N2971,N3038,N3079,N3546,N3671,N3803,N3804,N3809,N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,N146_O,N147_O,N148_O,N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,N156_O,N157_O,N158_O,N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,N166_O,N167_O,N168_O,N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,N176_O,N177_O,N178_O,N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,N186_O,N187_O,N188_O,N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,N196_O,N197_O,N198_O,N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,N206_O,N207_O,N208_O,N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,N216_O,N217_O,N218_O);

	initial begin
		#0.4 en = 0;
	end

	always #1 clk = ~clk;
	always #234 N1 = ~N1;
	always #233 N2 = ~N2;
	always #232 N3 = ~N3;
	always #231 N4 = ~N4;
	always #230 N5 = ~N5;
	always #229 N6 = ~N6;
	always #228 N7 = ~N7;
	always #227 N8 = ~N8;
	always #226 N11 = ~N11;
	always #225 N14 = ~N14;
	always #224 N15 = ~N15;
	always #223 N16 = ~N16;
	always #222 N19 = ~N19;
	always #221 N20 = ~N20;
	always #220 N21 = ~N21;
	always #219 N22 = ~N22;
	always #218 N23 = ~N23;
	always #217 N24 = ~N24;
	always #216 N25 = ~N25;
	always #215 N26 = ~N26;
	always #214 N27 = ~N27;
	always #213 N28 = ~N28;
	always #212 N29 = ~N29;
	always #211 N32 = ~N32;
	always #210 N33 = ~N33;
	always #209 N34 = ~N34;
	always #208 N35 = ~N35;
	always #207 N36 = ~N36;
	always #206 N37 = ~N37;
	always #205 N40 = ~N40;
	always #204 N43 = ~N43;
	always #203 N44 = ~N44;
	always #202 N47 = ~N47;
	always #201 N48 = ~N48;
	always #200 N49 = ~N49;
	always #199 N50 = ~N50;
	always #198 N51 = ~N51;
	always #197 N52 = ~N52;
	always #196 N53 = ~N53;
	always #195 N54 = ~N54;
	always #194 N55 = ~N55;
	always #193 N56 = ~N56;
	always #192 N57 = ~N57;
	always #191 N60 = ~N60;
	always #190 N61 = ~N61;
	always #189 N62 = ~N62;
	always #188 N63 = ~N63;
	always #187 N64 = ~N64;
	always #186 N65 = ~N65;
	always #185 N66 = ~N66;
	always #184 N67 = ~N67;
	always #183 N68 = ~N68;
	always #182 N69 = ~N69;
	always #181 N72 = ~N72;
	always #180 N73 = ~N73;
	always #179 N74 = ~N74;
	always #178 N75 = ~N75;
	always #177 N76 = ~N76;
	always #176 N77 = ~N77;
	always #175 N78 = ~N78;
	always #174 N79 = ~N79;
	always #173 N80 = ~N80;
	always #172 N81 = ~N81;
	always #171 N82 = ~N82;
	always #170 N85 = ~N85;
	always #169 N86 = ~N86;
	always #168 N87 = ~N87;
	always #167 N88 = ~N88;
	always #166 N89 = ~N89;
	always #165 N90 = ~N90;
	always #164 N91 = ~N91;
	always #163 N92 = ~N92;
	always #162 N93 = ~N93;
	always #161 N94 = ~N94;
	always #160 N95 = ~N95;
	always #159 N96 = ~N96;
	always #158 N99 = ~N99;
	always #157 N100 = ~N100;
	always #156 N101 = ~N101;
	always #155 N102 = ~N102;
	always #154 N103 = ~N103;
	always #153 N104 = ~N104;
	always #152 N105 = ~N105;
	always #151 N106 = ~N106;
	always #150 N107 = ~N107;
	always #149 N108 = ~N108;
	always #148 N111 = ~N111;
	always #147 N112 = ~N112;
	always #146 N113 = ~N113;
	always #145 N114 = ~N114;
	always #144 N115 = ~N115;
	always #143 N116 = ~N116;
	always #142 N117 = ~N117;
	always #141 N118 = ~N118;
	always #140 N119 = ~N119;
	always #139 N120 = ~N120;
	always #138 N123 = ~N123;
	always #137 N124 = ~N124;
	always #136 N125 = ~N125;
	always #135 N126 = ~N126;
	always #134 N127 = ~N127;
	always #133 N128 = ~N128;
	always #132 N129 = ~N129;
	always #131 N130 = ~N130;
	always #130 N131 = ~N131;
	always #129 N132 = ~N132;
	always #128 N135 = ~N135;
	always #127 N136 = ~N136;
	always #126 N137 = ~N137;
	always #125 N138 = ~N138;
	always #124 N139 = ~N139;
	always #123 N140 = ~N140;
	always #122 N141 = ~N141;
	always #121 N142 = ~N142;
	always #120 N219 = ~N219;
	always #119 N224 = ~N224;
	always #118 N227 = ~N227;
	always #117 N230 = ~N230;
	always #116 N231 = ~N231;
	always #115 N234 = ~N234;
	always #114 N237 = ~N237;
	always #113 N241 = ~N241;
	always #112 N246 = ~N246;
	always #111 N253 = ~N253;
	always #110 N256 = ~N256;
	always #109 N259 = ~N259;
	always #108 N262 = ~N262;
	always #107 N263 = ~N263;
	always #106 N266 = ~N266;
	always #105 N269 = ~N269;
	always #104 N272 = ~N272;
	always #103 N275 = ~N275;
	always #102 N278 = ~N278;
	always #101 N281 = ~N281;
	always #100 N284 = ~N284;
	always #99 N287 = ~N287;
	always #98 N290 = ~N290;
	always #97 N294 = ~N294;
	always #96 N297 = ~N297;
	always #95 N301 = ~N301;
	always #94 N305 = ~N305;
	always #93 N309 = ~N309;
	always #92 N313 = ~N313;
	always #91 N316 = ~N316;
	always #90 N319 = ~N319;
	always #89 N322 = ~N322;
	always #88 N325 = ~N325;
	always #87 N328 = ~N328;
	always #86 N331 = ~N331;
	always #85 N334 = ~N334;
	always #84 N337 = ~N337;
	always #83 N340 = ~N340;
	always #82 N343 = ~N343;
	always #81 N346 = ~N346;
	always #80 N349 = ~N349;
	always #79 N352 = ~N352;
	always #78 N355 = ~N355;
	always #77 N143_I = ~N143_I;
	always #76 N144_I = ~N144_I;
	always #75 N145_I = ~N145_I;
	always #74 N146_I = ~N146_I;
	always #73 N147_I = ~N147_I;
	always #72 N148_I = ~N148_I;
	always #71 N149_I = ~N149_I;
	always #70 N150_I = ~N150_I;
	always #69 N151_I = ~N151_I;
	always #68 N152_I = ~N152_I;
	always #67 N153_I = ~N153_I;
	always #66 N154_I = ~N154_I;
	always #65 N155_I = ~N155_I;
	always #64 N156_I = ~N156_I;
	always #63 N157_I = ~N157_I;
	always #62 N158_I = ~N158_I;
	always #61 N159_I = ~N159_I;
	always #60 N160_I = ~N160_I;
	always #59 N161_I = ~N161_I;
	always #58 N162_I = ~N162_I;
	always #57 N163_I = ~N163_I;
	always #56 N164_I = ~N164_I;
	always #55 N165_I = ~N165_I;
	always #54 N166_I = ~N166_I;
	always #53 N167_I = ~N167_I;
	always #52 N168_I = ~N168_I;
	always #51 N169_I = ~N169_I;
	always #50 N170_I = ~N170_I;
	always #49 N171_I = ~N171_I;
	always #48 N172_I = ~N172_I;
	always #47 N173_I = ~N173_I;
	always #46 N174_I = ~N174_I;
	always #45 N175_I = ~N175_I;
	always #44 N176_I = ~N176_I;
	always #43 N177_I = ~N177_I;
	always #42 N178_I = ~N178_I;
	always #41 N179_I = ~N179_I;
	always #40 N180_I = ~N180_I;
	always #39 N181_I = ~N181_I;
	always #38 N182_I = ~N182_I;
	always #37 N183_I = ~N183_I;
	always #36 N184_I = ~N184_I;
	always #35 N185_I = ~N185_I;
	always #34 N186_I = ~N186_I;
	always #33 N187_I = ~N187_I;
	always #32 N188_I = ~N188_I;
	always #31 N189_I = ~N189_I;
	always #30 N190_I = ~N190_I;
	always #29 N191_I = ~N191_I;
	always #28 N192_I = ~N192_I;
	always #27 N193_I = ~N193_I;
	always #26 N194_I = ~N194_I;
	always #25 N195_I = ~N195_I;
	always #24 N196_I = ~N196_I;
	always #23 N197_I = ~N197_I;
	always #22 N198_I = ~N198_I;
	always #21 N199_I = ~N199_I;
	always #20 N200_I = ~N200_I;
	always #19 N201_I = ~N201_I;
	always #18 N202_I = ~N202_I;
	always #17 N203_I = ~N203_I;
	always #16 N204_I = ~N204_I;
	always #15 N205_I = ~N205_I;
	always #14 N206_I = ~N206_I;
	always #13 N207_I = ~N207_I;
	always #12 N208_I = ~N208_I;
	always #11 N209_I = ~N209_I;
	always #10 N210_I = ~N210_I;
	always #9 N211_I = ~N211_I;
	always #8 N212_I = ~N212_I;
	always #7 N213_I = ~N213_I;
	always #6 N214_I = ~N214_I;
	always #5 N215_I = ~N215_I;
	always #4 N216_I = ~N216_I;
	always #3 N217_I = ~N217_I;
	always #2 N218_I = ~N218_I;	

	initial #1024 $finish;
endmodule